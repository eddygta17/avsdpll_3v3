magic
tech scmos
timestamp 1599458516
<< nwell >>
rect 0 51 231 108
rect 0 -167 231 -54
<< ntransistor >>
rect 16 9 18 19
rect 50 9 52 29
rect 55 9 57 29
rect 91 9 93 19
rect 126 9 128 19
rect 163 9 165 39
rect 168 9 170 39
rect 173 9 175 39
rect 212 9 214 19
rect 17 -32 19 -12
rect 22 -32 24 -12
rect 41 -32 43 -12
rect 46 -32 48 -12
rect 65 -32 67 -12
rect 70 -32 72 -12
rect 78 -22 80 -12
rect 97 -32 99 -12
rect 102 -32 104 -12
rect 110 -22 112 -12
rect 129 -32 131 -12
rect 134 -32 136 -12
rect 142 -22 144 -12
rect 161 -22 163 -12
rect 178 -32 180 -12
rect 183 -32 185 -12
rect 202 -32 204 -12
rect 207 -32 209 -12
rect 16 -209 18 -199
rect 50 -209 52 -189
rect 55 -209 57 -189
rect 91 -209 93 -199
rect 126 -209 128 -199
rect 163 -209 165 -179
rect 168 -209 170 -179
rect 173 -209 175 -179
rect 212 -209 214 -199
<< ptransistor >>
rect 16 77 18 97
rect 50 77 52 97
rect 58 77 60 97
rect 91 77 93 97
rect 126 77 128 97
rect 163 77 165 97
rect 171 77 173 97
rect 179 77 181 97
rect 212 77 214 97
rect 17 -100 19 -80
rect 25 -100 27 -80
rect 41 -100 43 -80
rect 49 -100 51 -80
rect 65 -100 67 -80
rect 73 -100 75 -80
rect 81 -100 83 -80
rect 97 -100 99 -80
rect 105 -100 107 -80
rect 113 -100 115 -80
rect 129 -100 131 -80
rect 137 -100 139 -80
rect 145 -100 147 -80
rect 161 -100 163 -80
rect 178 -100 180 -80
rect 186 -100 188 -80
rect 202 -100 204 -80
rect 210 -100 212 -80
rect 16 -141 18 -121
rect 50 -141 52 -121
rect 58 -141 60 -121
rect 91 -141 93 -121
rect 126 -141 128 -121
rect 163 -141 165 -121
rect 171 -141 173 -121
rect 179 -141 181 -121
rect 212 -141 214 -121
<< ndiffusion >>
rect 11 18 16 19
rect 15 9 16 18
rect 18 18 23 19
rect 18 9 19 18
rect 49 9 50 29
rect 52 9 55 29
rect 57 9 58 29
rect 86 18 91 19
rect 90 9 91 18
rect 93 18 98 19
rect 93 9 94 18
rect 121 18 126 19
rect 125 9 126 18
rect 128 18 133 19
rect 128 9 129 18
rect 162 9 163 39
rect 165 9 168 39
rect 170 9 173 39
rect 175 9 176 39
rect 207 18 212 19
rect 211 9 212 18
rect 214 18 219 19
rect 214 9 215 18
rect 16 -32 17 -12
rect 19 -32 22 -12
rect 24 -32 25 -12
rect 40 -32 41 -12
rect 43 -32 46 -12
rect 48 -32 49 -12
rect 64 -32 65 -12
rect 67 -32 70 -12
rect 72 -32 73 -12
rect 77 -22 78 -12
rect 80 -22 81 -12
rect 96 -32 97 -12
rect 99 -32 102 -12
rect 104 -32 105 -12
rect 109 -22 110 -12
rect 112 -22 113 -12
rect 128 -32 129 -12
rect 131 -32 134 -12
rect 136 -32 137 -12
rect 141 -22 142 -12
rect 144 -22 145 -12
rect 160 -21 161 -12
rect 156 -22 161 -21
rect 163 -21 164 -12
rect 163 -22 168 -21
rect 177 -32 178 -12
rect 180 -32 183 -12
rect 185 -32 186 -12
rect 201 -32 202 -12
rect 204 -32 207 -12
rect 209 -32 210 -12
rect 11 -200 16 -199
rect 15 -209 16 -200
rect 18 -200 23 -199
rect 18 -209 19 -200
rect 49 -209 50 -189
rect 52 -209 55 -189
rect 57 -209 58 -189
rect 86 -200 91 -199
rect 90 -209 91 -200
rect 93 -200 98 -199
rect 93 -209 94 -200
rect 121 -200 126 -199
rect 125 -209 126 -200
rect 128 -200 133 -199
rect 128 -209 129 -200
rect 162 -209 163 -179
rect 165 -209 168 -179
rect 170 -209 173 -179
rect 175 -209 176 -179
rect 207 -200 212 -199
rect 211 -209 212 -200
rect 214 -200 219 -199
rect 214 -209 215 -200
<< pdiffusion >>
rect 11 96 16 97
rect 15 77 16 96
rect 18 96 23 97
rect 18 77 19 96
rect 49 77 50 97
rect 52 77 53 97
rect 57 77 58 97
rect 60 77 61 97
rect 86 96 91 97
rect 90 77 91 96
rect 93 96 98 97
rect 93 77 94 96
rect 121 96 126 97
rect 125 77 126 96
rect 128 96 133 97
rect 128 77 129 96
rect 162 77 163 97
rect 165 77 166 97
rect 170 77 171 97
rect 173 79 174 97
rect 178 79 179 97
rect 173 77 179 79
rect 181 77 182 97
rect 207 96 212 97
rect 211 77 212 96
rect 214 96 219 97
rect 214 77 215 96
rect 16 -100 17 -80
rect 19 -100 20 -80
rect 24 -100 25 -80
rect 27 -100 28 -80
rect 40 -100 41 -80
rect 43 -100 44 -80
rect 48 -100 49 -80
rect 51 -100 52 -80
rect 64 -100 65 -80
rect 67 -100 68 -80
rect 72 -100 73 -80
rect 75 -100 76 -80
rect 80 -100 81 -80
rect 83 -100 84 -80
rect 96 -100 97 -80
rect 99 -100 100 -80
rect 104 -100 105 -80
rect 107 -100 108 -80
rect 112 -100 113 -80
rect 115 -100 116 -80
rect 128 -100 129 -80
rect 131 -100 132 -80
rect 136 -100 137 -80
rect 139 -100 140 -80
rect 144 -100 145 -80
rect 147 -100 148 -80
rect 160 -99 161 -80
rect 156 -100 161 -99
rect 163 -99 164 -80
rect 163 -100 168 -99
rect 177 -100 178 -80
rect 180 -100 181 -80
rect 185 -100 186 -80
rect 188 -100 189 -80
rect 201 -100 202 -80
rect 204 -100 205 -80
rect 209 -100 210 -80
rect 212 -100 213 -80
rect 11 -122 16 -121
rect 15 -141 16 -122
rect 18 -122 23 -121
rect 18 -141 19 -122
rect 49 -141 50 -121
rect 52 -141 53 -121
rect 57 -141 58 -121
rect 60 -141 61 -121
rect 86 -122 91 -121
rect 90 -141 91 -122
rect 93 -122 98 -121
rect 93 -141 94 -122
rect 121 -122 126 -121
rect 125 -141 126 -122
rect 128 -122 133 -121
rect 128 -141 129 -122
rect 162 -141 163 -121
rect 165 -141 166 -121
rect 170 -141 171 -121
rect 173 -139 174 -121
rect 178 -139 179 -121
rect 173 -141 179 -139
rect 181 -141 182 -121
rect 207 -122 212 -121
rect 211 -141 212 -122
rect 214 -122 219 -121
rect 214 -141 215 -122
<< ndcontact >>
rect 11 9 15 18
rect 19 9 23 18
rect 45 9 49 29
rect 58 9 62 29
rect 86 9 90 18
rect 94 9 98 18
rect 121 9 125 18
rect 129 9 133 18
rect 158 9 162 39
rect 176 9 180 39
rect 207 9 211 18
rect 215 9 219 18
rect 12 -32 16 -12
rect 25 -32 29 -12
rect 36 -32 40 -12
rect 49 -32 53 -12
rect 60 -32 64 -12
rect 73 -32 77 -12
rect 81 -22 85 -12
rect 92 -32 96 -12
rect 105 -32 109 -12
rect 113 -22 117 -12
rect 124 -32 128 -12
rect 137 -32 141 -12
rect 145 -22 149 -12
rect 156 -21 160 -12
rect 164 -21 168 -12
rect 173 -32 177 -12
rect 186 -32 190 -12
rect 197 -32 201 -12
rect 210 -32 214 -12
rect 11 -209 15 -200
rect 19 -209 23 -200
rect 45 -209 49 -189
rect 58 -209 62 -189
rect 86 -209 90 -200
rect 94 -209 98 -200
rect 121 -209 125 -200
rect 129 -209 133 -200
rect 158 -209 162 -179
rect 176 -209 180 -179
rect 207 -209 211 -200
rect 215 -209 219 -200
<< pdcontact >>
rect 11 77 15 96
rect 19 77 23 96
rect 45 77 49 97
rect 53 77 57 97
rect 61 77 65 97
rect 86 77 90 96
rect 94 77 98 96
rect 121 77 125 96
rect 129 77 133 96
rect 158 77 162 97
rect 166 77 170 97
rect 174 79 178 97
rect 182 77 186 97
rect 207 77 211 96
rect 215 77 219 96
rect 12 -100 16 -80
rect 20 -100 24 -80
rect 28 -100 32 -80
rect 36 -100 40 -80
rect 44 -100 48 -80
rect 52 -100 56 -80
rect 60 -100 64 -80
rect 68 -100 72 -80
rect 76 -100 80 -80
rect 84 -100 88 -80
rect 92 -100 96 -80
rect 100 -100 104 -80
rect 108 -100 112 -80
rect 116 -100 120 -80
rect 124 -100 128 -80
rect 132 -100 136 -80
rect 140 -100 144 -80
rect 148 -100 152 -80
rect 156 -99 160 -80
rect 164 -99 168 -80
rect 173 -100 177 -80
rect 181 -100 185 -80
rect 189 -100 193 -80
rect 197 -100 201 -80
rect 205 -100 209 -80
rect 213 -100 217 -80
rect 11 -141 15 -122
rect 19 -141 23 -122
rect 45 -141 49 -121
rect 53 -141 57 -121
rect 61 -141 65 -121
rect 86 -141 90 -122
rect 94 -141 98 -122
rect 121 -141 125 -122
rect 129 -141 133 -122
rect 158 -141 162 -121
rect 166 -141 170 -121
rect 174 -139 178 -121
rect 182 -141 186 -121
rect 207 -141 211 -122
rect 215 -141 219 -122
<< psubstratepcontact >>
rect 7 1 11 5
rect 41 1 45 5
rect 57 1 61 5
rect 82 1 86 5
rect 117 1 121 5
rect 154 1 158 5
rect 170 1 174 5
rect 205 1 209 5
rect 8 -8 12 -4
rect 24 -8 28 -4
rect 32 -8 36 -4
rect 48 -8 52 -4
rect 72 -8 76 -4
rect 87 -8 91 -4
rect 104 -8 108 -4
rect 136 -8 140 -4
rect 152 -8 156 -4
rect 185 -8 189 -4
rect 193 -8 197 -4
rect 209 -8 213 -4
rect 7 -217 11 -213
rect 41 -217 45 -213
rect 57 -217 61 -213
rect 82 -217 86 -213
rect 117 -217 121 -213
rect 154 -217 158 -213
rect 170 -217 174 -213
rect 205 -217 209 -213
<< nsubstratencontact >>
rect 7 101 11 105
rect 41 101 45 105
rect 57 101 61 105
rect 82 101 86 105
rect 117 101 121 105
rect 154 101 158 105
rect 170 101 174 105
rect 203 101 207 105
rect 8 -108 12 -104
rect 24 -108 28 -104
rect 32 -108 36 -104
rect 48 -108 52 -104
rect 72 -108 76 -104
rect 87 -108 91 -104
rect 104 -108 108 -104
rect 117 -108 124 -104
rect 136 -108 140 -104
rect 152 -108 156 -104
rect 185 -108 189 -104
rect 193 -108 197 -104
rect 209 -108 213 -104
rect 7 -117 11 -113
rect 41 -117 45 -113
rect 57 -117 61 -113
rect 82 -117 86 -113
rect 117 -117 121 -113
rect 154 -117 158 -113
rect 170 -117 174 -113
rect 203 -117 207 -113
<< polysilicon >>
rect 16 97 18 99
rect 50 97 52 99
rect 58 97 60 99
rect 91 97 93 99
rect 126 97 128 99
rect 163 97 165 99
rect 171 97 173 99
rect 179 97 181 99
rect 212 97 214 99
rect 16 26 18 77
rect 50 36 52 77
rect 49 32 52 36
rect 58 64 60 77
rect 58 60 61 64
rect 58 32 60 60
rect 50 29 52 32
rect 55 30 60 32
rect 55 29 57 30
rect 15 22 18 26
rect 16 19 18 22
rect 91 26 93 77
rect 126 26 128 77
rect 163 56 165 77
rect 171 76 173 77
rect 162 52 165 56
rect 163 39 165 52
rect 168 74 173 76
rect 168 39 170 74
rect 179 66 181 77
rect 178 62 181 66
rect 179 42 181 62
rect 173 40 181 42
rect 173 39 175 40
rect 90 22 93 26
rect 125 22 128 26
rect 91 19 93 22
rect 126 19 128 22
rect 212 26 214 77
rect 211 22 214 26
rect 212 19 214 22
rect 16 7 18 9
rect 50 7 52 9
rect 55 7 57 9
rect 91 7 93 9
rect 126 7 128 9
rect 163 7 165 9
rect 168 7 170 9
rect 173 7 175 9
rect 212 7 214 9
rect 17 -12 19 -10
rect 22 -12 24 -10
rect 41 -12 43 -10
rect 46 -12 48 -10
rect 65 -12 67 -10
rect 70 -12 72 -10
rect 78 -12 80 -10
rect 97 -12 99 -10
rect 102 -12 104 -10
rect 110 -12 112 -10
rect 129 -12 131 -10
rect 134 -12 136 -10
rect 142 -12 144 -10
rect 161 -12 163 -10
rect 178 -12 180 -10
rect 183 -12 185 -10
rect 202 -12 204 -10
rect 207 -12 209 -10
rect 17 -35 19 -32
rect 22 -33 24 -32
rect 22 -35 27 -33
rect 41 -35 43 -32
rect 46 -33 48 -32
rect 46 -35 51 -33
rect 16 -39 19 -35
rect 17 -80 19 -39
rect 25 -63 27 -35
rect 40 -39 43 -35
rect 25 -67 28 -63
rect 25 -80 27 -67
rect 41 -80 43 -39
rect 49 -63 51 -35
rect 65 -40 67 -32
rect 64 -44 67 -40
rect 49 -67 52 -63
rect 49 -80 51 -67
rect 65 -80 67 -44
rect 70 -43 72 -32
rect 78 -35 80 -22
rect 82 -39 83 -36
rect 70 -45 75 -43
rect 73 -48 75 -45
rect 73 -80 75 -52
rect 81 -80 83 -39
rect 97 -47 99 -32
rect 102 -43 104 -32
rect 110 -35 112 -22
rect 114 -39 115 -36
rect 102 -45 107 -43
rect 96 -51 99 -47
rect 97 -80 99 -51
rect 105 -55 107 -45
rect 105 -80 107 -59
rect 113 -80 115 -39
rect 129 -43 131 -32
rect 128 -47 131 -43
rect 134 -43 136 -32
rect 142 -35 144 -22
rect 161 -25 163 -22
rect 160 -29 163 -25
rect 146 -39 147 -36
rect 134 -45 139 -43
rect 129 -80 131 -47
rect 137 -55 139 -45
rect 137 -80 139 -59
rect 145 -80 147 -39
rect 161 -80 163 -29
rect 178 -35 180 -32
rect 183 -33 185 -32
rect 183 -35 188 -33
rect 202 -35 204 -32
rect 207 -33 209 -32
rect 207 -35 212 -33
rect 177 -39 180 -35
rect 178 -80 180 -39
rect 186 -69 188 -35
rect 201 -39 204 -35
rect 186 -73 189 -69
rect 186 -80 188 -73
rect 202 -80 204 -39
rect 210 -58 212 -35
rect 210 -62 213 -58
rect 210 -80 212 -62
rect 17 -102 19 -100
rect 25 -102 27 -100
rect 41 -102 43 -100
rect 49 -102 51 -100
rect 65 -102 67 -100
rect 73 -102 75 -100
rect 81 -102 83 -100
rect 97 -102 99 -100
rect 105 -102 107 -100
rect 113 -102 115 -100
rect 129 -102 131 -100
rect 137 -102 139 -100
rect 145 -102 147 -100
rect 161 -102 163 -100
rect 178 -102 180 -100
rect 186 -102 188 -100
rect 202 -102 204 -100
rect 210 -102 212 -100
rect 16 -121 18 -119
rect 50 -121 52 -119
rect 58 -121 60 -119
rect 91 -121 93 -119
rect 126 -121 128 -119
rect 163 -121 165 -119
rect 171 -121 173 -119
rect 179 -121 181 -119
rect 212 -121 214 -119
rect 16 -192 18 -141
rect 50 -182 52 -141
rect 49 -186 52 -182
rect 58 -154 60 -141
rect 58 -158 61 -154
rect 58 -186 60 -158
rect 50 -189 52 -186
rect 55 -188 60 -186
rect 55 -189 57 -188
rect 15 -196 18 -192
rect 16 -199 18 -196
rect 91 -192 93 -141
rect 126 -192 128 -141
rect 163 -162 165 -141
rect 171 -142 173 -141
rect 162 -166 165 -162
rect 163 -179 165 -166
rect 168 -144 173 -142
rect 168 -179 170 -144
rect 179 -152 181 -141
rect 178 -156 181 -152
rect 179 -176 181 -156
rect 173 -178 181 -176
rect 173 -179 175 -178
rect 90 -196 93 -192
rect 125 -196 128 -192
rect 91 -199 93 -196
rect 126 -199 128 -196
rect 212 -192 214 -141
rect 211 -196 214 -192
rect 212 -199 214 -196
rect 16 -211 18 -209
rect 50 -211 52 -209
rect 55 -211 57 -209
rect 91 -211 93 -209
rect 126 -211 128 -209
rect 163 -211 165 -209
rect 168 -211 170 -209
rect 173 -211 175 -209
rect 212 -211 214 -209
<< polycontact >>
rect 45 32 49 36
rect 61 60 65 64
rect 11 22 15 26
rect 158 52 162 56
rect 174 62 178 66
rect 170 46 174 50
rect 86 22 90 26
rect 121 22 125 26
rect 207 22 211 26
rect 12 -39 16 -35
rect 36 -39 40 -35
rect 28 -67 32 -63
rect 60 -44 64 -40
rect 52 -67 56 -63
rect 78 -39 82 -35
rect 71 -52 75 -48
rect 110 -39 114 -35
rect 92 -51 96 -47
rect 103 -59 107 -55
rect 124 -47 128 -43
rect 156 -29 160 -25
rect 142 -39 146 -35
rect 135 -59 139 -55
rect 173 -39 177 -35
rect 197 -39 201 -35
rect 189 -73 193 -69
rect 213 -62 217 -58
rect 45 -186 49 -182
rect 61 -158 65 -154
rect 11 -196 15 -192
rect 158 -166 162 -162
rect 174 -156 178 -152
rect 170 -172 174 -168
rect 86 -196 90 -192
rect 121 -196 125 -192
rect 207 -196 211 -192
<< metal1 >>
rect 7 105 223 106
rect 11 101 41 105
rect 45 101 57 105
rect 61 101 82 105
rect 86 101 117 105
rect 121 101 154 105
rect 158 101 170 105
rect 174 101 203 105
rect 207 101 223 105
rect 7 100 223 101
rect 11 96 15 100
rect 45 97 49 100
rect 61 97 65 100
rect 19 96 23 97
rect 86 96 90 100
rect 94 96 98 97
rect 121 96 125 100
rect 158 97 162 100
rect 174 97 178 100
rect 129 96 133 97
rect 19 36 23 77
rect 53 74 57 77
rect 19 32 45 36
rect 0 22 11 26
rect 11 18 15 19
rect 19 18 23 32
rect 53 30 57 70
rect 61 56 65 60
rect 94 30 98 77
rect 129 70 133 77
rect 167 76 170 77
rect 207 96 211 100
rect 215 96 219 97
rect 182 76 185 77
rect 167 73 185 76
rect 129 66 178 70
rect 53 29 90 30
rect 53 26 58 29
rect 62 26 90 29
rect 94 26 125 30
rect 86 18 90 19
rect 94 18 98 26
rect 121 18 125 19
rect 129 18 133 66
rect 182 64 185 73
rect 158 56 162 60
rect 182 56 186 60
rect 167 46 170 50
rect 182 40 185 56
rect 177 39 185 40
rect 180 37 185 39
rect 180 26 195 30
rect 199 26 211 30
rect 215 26 219 77
rect 215 22 231 26
rect 207 18 211 19
rect 215 18 219 22
rect 11 6 15 9
rect 45 6 49 9
rect 86 6 90 9
rect 121 6 125 9
rect 158 6 162 9
rect 207 6 211 9
rect 7 5 223 6
rect 11 1 41 5
rect 45 1 57 5
rect 61 1 82 5
rect 86 1 117 5
rect 121 1 154 5
rect 158 1 170 5
rect 174 1 205 5
rect 209 1 223 5
rect 7 -4 223 1
rect 7 -8 8 -4
rect 12 -8 24 -4
rect 28 -8 32 -4
rect 36 -8 48 -4
rect 52 -8 72 -4
rect 76 -8 87 -4
rect 91 -8 104 -4
rect 108 -8 136 -4
rect 140 -8 152 -4
rect 156 -8 185 -4
rect 189 -8 193 -4
rect 197 -8 209 -4
rect 213 -8 223 -4
rect 7 -9 223 -8
rect 12 -12 16 -9
rect 36 -12 40 -9
rect 73 -12 77 -9
rect 105 -12 109 -9
rect 137 -12 141 -9
rect 156 -12 160 -9
rect 173 -12 177 -9
rect 197 -12 201 -9
rect 20 -32 25 -29
rect 44 -32 49 -29
rect 81 -25 88 -22
rect 12 -43 16 -39
rect 20 -39 24 -32
rect 20 -43 40 -39
rect 20 -48 24 -43
rect 20 -80 24 -52
rect 44 -59 48 -32
rect 61 -35 70 -32
rect 67 -36 70 -35
rect 67 -39 78 -36
rect 60 -40 64 -39
rect 70 -52 71 -48
rect 28 -63 48 -59
rect 44 -80 48 -63
rect 52 -63 56 -59
rect 78 -74 81 -39
rect 85 -51 88 -25
rect 113 -25 120 -22
rect 93 -35 102 -32
rect 99 -36 102 -35
rect 99 -39 110 -36
rect 117 -39 120 -25
rect 156 -22 160 -21
rect 145 -25 152 -22
rect 149 -29 152 -25
rect 125 -35 134 -32
rect 149 -33 160 -29
rect 131 -36 134 -35
rect 131 -39 142 -36
rect 92 -47 96 -43
rect 85 -69 88 -55
rect 100 -63 107 -59
rect 84 -73 88 -69
rect 69 -77 81 -74
rect 69 -80 72 -77
rect 85 -80 88 -73
rect 110 -74 113 -39
rect 117 -43 128 -39
rect 117 -69 120 -43
rect 132 -63 139 -59
rect 116 -73 120 -69
rect 101 -77 113 -74
rect 101 -80 104 -77
rect 117 -80 120 -73
rect 142 -74 145 -39
rect 149 -69 152 -33
rect 148 -73 152 -69
rect 133 -77 145 -74
rect 133 -80 136 -77
rect 149 -80 152 -73
rect 164 -39 168 -21
rect 181 -32 186 -29
rect 205 -32 210 -29
rect 173 -43 177 -39
rect 181 -39 185 -32
rect 181 -43 201 -39
rect 164 -80 168 -43
rect 181 -80 185 -43
rect 205 -73 209 -32
rect 213 -58 217 -54
rect 189 -77 209 -73
rect 205 -80 209 -77
rect 12 -103 16 -100
rect 28 -103 32 -100
rect 36 -103 40 -100
rect 52 -103 56 -100
rect 60 -103 64 -100
rect 76 -103 80 -100
rect 92 -103 96 -100
rect 108 -103 112 -100
rect 124 -103 128 -100
rect 140 -103 144 -100
rect 156 -103 160 -99
rect 164 -100 168 -99
rect 173 -103 177 -100
rect 189 -103 193 -100
rect 197 -103 201 -100
rect 213 -103 217 -100
rect 7 -104 223 -103
rect 7 -108 8 -104
rect 12 -108 24 -104
rect 28 -108 32 -104
rect 36 -108 48 -104
rect 52 -108 72 -104
rect 76 -108 87 -104
rect 91 -108 104 -104
rect 108 -108 117 -104
rect 124 -108 136 -104
rect 140 -108 152 -104
rect 156 -108 185 -104
rect 189 -108 193 -104
rect 197 -108 209 -104
rect 213 -108 223 -104
rect 7 -113 223 -108
rect 11 -117 41 -113
rect 45 -117 57 -113
rect 61 -117 82 -113
rect 86 -117 117 -113
rect 121 -117 154 -113
rect 158 -117 170 -113
rect 174 -117 203 -113
rect 207 -117 223 -113
rect 7 -118 223 -117
rect 11 -122 15 -118
rect 45 -121 49 -118
rect 61 -121 65 -118
rect 19 -122 23 -121
rect 86 -122 90 -118
rect 94 -122 98 -121
rect 121 -122 125 -118
rect 158 -121 162 -118
rect 174 -121 178 -118
rect 129 -122 133 -121
rect 19 -182 23 -141
rect 53 -145 57 -141
rect 19 -186 45 -182
rect 0 -196 11 -192
rect 11 -200 15 -199
rect 19 -200 23 -186
rect 53 -188 57 -149
rect 61 -162 65 -158
rect 94 -188 98 -141
rect 129 -148 133 -141
rect 167 -142 170 -141
rect 207 -122 211 -118
rect 215 -122 219 -121
rect 182 -142 185 -141
rect 167 -145 185 -142
rect 129 -152 178 -148
rect 53 -189 90 -188
rect 53 -192 58 -189
rect 62 -192 90 -189
rect 94 -192 125 -188
rect 86 -200 90 -199
rect 94 -200 98 -192
rect 121 -200 125 -199
rect 129 -200 133 -152
rect 182 -158 185 -145
rect 158 -162 162 -158
rect 182 -162 186 -158
rect 166 -172 170 -168
rect 182 -178 185 -162
rect 177 -179 185 -178
rect 180 -181 185 -179
rect 180 -192 188 -188
rect 192 -192 211 -188
rect 215 -192 219 -141
rect 215 -196 231 -192
rect 207 -200 211 -199
rect 215 -200 219 -196
rect 11 -212 15 -209
rect 45 -212 49 -209
rect 86 -212 90 -209
rect 121 -212 125 -209
rect 158 -212 162 -209
rect 207 -212 211 -209
rect 7 -213 223 -212
rect 11 -217 41 -213
rect 45 -217 57 -213
rect 61 -217 82 -213
rect 86 -217 117 -213
rect 121 -217 154 -213
rect 158 -217 170 -213
rect 174 -217 205 -213
rect 209 -217 223 -213
rect 7 -218 223 -217
<< m2contact >>
rect 53 70 57 74
rect 61 60 65 64
rect 158 52 162 56
rect 170 46 174 50
rect 195 26 199 30
rect 12 -39 16 -35
rect 20 -52 24 -48
rect 60 -44 64 -40
rect 71 -52 75 -48
rect 52 -67 56 -63
rect 110 -39 114 -35
rect 92 -51 96 -47
rect 85 -55 89 -51
rect 135 -59 139 -55
rect 164 -43 168 -39
rect 173 -39 177 -35
rect 189 -73 193 -69
rect 213 -62 217 -58
rect 53 -149 57 -145
rect 61 -158 65 -154
rect 158 -166 162 -162
rect 170 -172 174 -168
rect 188 -192 192 -188
<< metal2 >>
rect 57 70 217 74
rect 65 60 199 64
rect 109 -39 110 -35
rect 158 -39 162 52
rect 169 46 170 50
rect 195 30 199 60
rect 12 -40 16 -39
rect 12 -44 60 -40
rect 158 -43 164 -39
rect 168 -43 177 -39
rect 12 -144 16 -44
rect 92 -47 96 -46
rect 24 -52 71 -48
rect 89 -55 139 -51
rect 158 -63 162 -43
rect 213 -58 217 70
rect 56 -67 162 -63
rect 12 -149 53 -144
rect 61 -198 65 -158
rect 158 -162 162 -67
rect 189 -74 193 -73
rect 80 -172 170 -168
rect 188 -198 192 -192
rect 61 -202 192 -198
<< m3contact >>
rect 110 -39 114 -35
rect 170 46 174 50
rect 71 -52 75 -48
rect 92 -51 96 -47
rect 213 -62 217 -58
rect 189 -73 193 -69
rect 76 -172 80 -168
<< metal3 >>
rect 92 46 170 50
rect 92 -47 96 46
rect 75 -52 80 -48
rect 76 -168 80 -52
rect 92 -69 96 -51
rect 110 -58 114 -39
rect 110 -62 213 -58
rect 92 -73 189 -69
<< m1p >>
rect 174 66 178 70
rect 61 56 65 60
rect 158 56 162 60
rect 182 56 186 60
rect 53 46 57 50
rect 167 46 171 50
rect 19 36 23 40
rect 94 36 98 40
rect 129 36 133 40
rect 215 36 219 40
rect 67 26 71 30
rect 0 22 15 26
rect 156 -33 160 -29
rect 12 -43 16 -39
rect 22 -43 40 -39
rect 60 -43 64 -39
rect 124 -43 128 -39
rect 164 -43 168 -39
rect 173 -43 177 -39
rect 183 -43 201 -39
rect 92 -47 96 -43
rect 20 -53 24 -49
rect 44 -53 48 -49
rect 70 -52 74 -48
rect 181 -53 185 -49
rect 205 -53 209 -49
rect 28 -63 32 -59
rect 52 -63 56 -59
rect 100 -63 104 -59
rect 132 -63 136 -59
rect 84 -73 88 -69
rect 116 -73 120 -69
rect 148 -73 152 -69
rect 174 -152 178 -148
rect 61 -162 65 -158
rect 158 -162 162 -158
rect 182 -162 186 -158
rect 53 -172 57 -168
rect 166 -172 170 -168
rect 19 -182 23 -178
rect 94 -182 98 -178
rect 129 -182 133 -178
rect 215 -182 219 -178
rect 67 -192 71 -188
rect 0 -196 15 -192
<< labels >>
rlabel metal1 0 22 0 26 3 clockin
rlabel metal1 0 -196 0 -192 3 vcoin
rlabel metal1 166 -50 166 -50 1 RESET
rlabel metal1 79 27 79 27 1 B
rlabel metal1 78 -190 78 -190 1 C
rlabel metal1 13 -41 13 -41 1 C
rlabel metal1 174 -42 174 -42 1 RESET
rlabel metal1 207 -62 207 -62 1 A
rlabel metal1 22 -58 22 -58 1 D
rlabel metal1 54 -61 54 -61 1 RESET
rlabel metal1 160 59 160 59 1 RESET
rlabel metal1 160 -161 160 -161 1 RESET
rlabel metal1 168 48 168 48 1 A
rlabel polycontact 126 -45 126 -45 1 A1
rlabel polycontact 137 -57 137 -57 1 A2
rlabel metal1 168 -170 168 -170 1 D
rlabel metal1 231 -196 231 -192 7 down
rlabel polycontact 73 -51 73 -51 1 D
rlabel polycontact 61 -42 61 -42 1 C
rlabel polycontact 112 -37 112 -37 1 B
rlabel polycontact 94 -49 94 -49 1 A
rlabel metal1 216 -56 216 -56 1 B
<< end >>
