magic
tech scmos
timestamp 1599387492
<< nwell >>
rect -134 -3 235 27
<< ntransistor >>
rect -125 -15 -122 -9
rect -101 -15 -98 -9
rect -77 -15 -74 -9
rect -53 -15 -50 -9
rect -29 -15 -26 -9
rect -2 -15 1 -9
rect 22 -15 25 -9
rect 46 -15 49 -9
rect 70 -15 73 -9
rect 94 -15 97 -9
rect 121 -15 124 -9
rect 145 -15 148 -9
rect 169 -15 172 -9
rect 193 -15 196 -9
rect 217 -15 220 -9
<< ptransistor >>
rect -101 3 -98 11
rect -77 3 -74 11
rect -53 3 -50 11
rect -29 3 -26 11
rect 22 3 25 11
rect 46 3 49 11
rect 70 3 73 11
rect 94 3 97 11
rect 145 3 148 11
rect 169 3 172 11
rect 193 3 196 11
rect 217 3 220 11
<< ndiffusion >>
rect -134 -10 -125 -9
rect -134 -14 -133 -10
rect -129 -14 -125 -10
rect -134 -15 -125 -14
rect -122 -15 -101 -9
rect -98 -10 -89 -9
rect -98 -14 -94 -10
rect -90 -14 -89 -10
rect -98 -15 -89 -14
rect -86 -10 -77 -9
rect -86 -14 -85 -10
rect -81 -14 -77 -10
rect -86 -15 -77 -14
rect -74 -15 -53 -9
rect -50 -10 -41 -9
rect -50 -14 -46 -10
rect -42 -14 -41 -10
rect -50 -15 -41 -14
rect -38 -10 -29 -9
rect -38 -14 -37 -10
rect -33 -14 -29 -10
rect -38 -15 -29 -14
rect -26 -10 -17 -9
rect -26 -14 -22 -10
rect -18 -14 -17 -10
rect -26 -15 -17 -14
rect -11 -10 -2 -9
rect -11 -14 -10 -10
rect -6 -14 -2 -10
rect -11 -15 -2 -14
rect 1 -15 22 -9
rect 25 -10 34 -9
rect 25 -14 29 -10
rect 33 -14 34 -10
rect 25 -15 34 -14
rect 37 -10 46 -9
rect 37 -14 38 -10
rect 42 -14 46 -10
rect 37 -15 46 -14
rect 49 -15 70 -9
rect 73 -10 82 -9
rect 73 -14 77 -10
rect 81 -14 82 -10
rect 73 -15 82 -14
rect 85 -10 94 -9
rect 85 -14 86 -10
rect 90 -14 94 -10
rect 85 -15 94 -14
rect 97 -10 106 -9
rect 97 -14 101 -10
rect 105 -14 106 -10
rect 97 -15 106 -14
rect 112 -10 121 -9
rect 112 -14 113 -10
rect 117 -14 121 -10
rect 112 -15 121 -14
rect 124 -15 145 -9
rect 148 -10 157 -9
rect 148 -14 152 -10
rect 156 -14 157 -10
rect 148 -15 157 -14
rect 160 -10 169 -9
rect 160 -14 161 -10
rect 165 -14 169 -10
rect 160 -15 169 -14
rect 172 -15 193 -9
rect 196 -10 205 -9
rect 196 -14 200 -10
rect 204 -14 205 -10
rect 196 -15 205 -14
rect 208 -10 217 -9
rect 208 -14 209 -10
rect 213 -14 217 -10
rect 208 -15 217 -14
rect 220 -10 229 -9
rect 220 -14 224 -10
rect 228 -14 229 -10
rect 220 -15 229 -14
<< pdiffusion >>
rect -110 8 -101 11
rect -110 4 -109 8
rect -105 4 -101 8
rect -110 3 -101 4
rect -98 10 -89 11
rect -98 6 -94 10
rect -90 6 -89 10
rect -98 3 -89 6
rect -86 10 -77 11
rect -86 6 -85 10
rect -81 6 -77 10
rect -86 3 -77 6
rect -74 8 -65 11
rect -74 4 -70 8
rect -66 4 -65 8
rect -74 3 -65 4
rect -62 10 -53 11
rect -62 6 -61 10
rect -57 6 -53 10
rect -62 3 -53 6
rect -50 3 -29 11
rect -26 10 -17 11
rect -26 6 -22 10
rect -18 6 -17 10
rect -26 3 -17 6
rect 13 8 22 11
rect 13 4 14 8
rect 18 4 22 8
rect 13 3 22 4
rect 25 10 34 11
rect 25 6 29 10
rect 33 6 34 10
rect 25 3 34 6
rect 37 10 46 11
rect 37 6 38 10
rect 42 6 46 10
rect 37 3 46 6
rect 49 8 58 11
rect 49 4 53 8
rect 57 4 58 8
rect 49 3 58 4
rect 61 10 70 11
rect 61 6 62 10
rect 66 6 70 10
rect 61 3 70 6
rect 73 3 94 11
rect 97 10 106 11
rect 97 6 101 10
rect 105 6 106 10
rect 97 3 106 6
rect 136 8 145 11
rect 136 4 137 8
rect 141 4 145 8
rect 136 3 145 4
rect 148 10 157 11
rect 148 6 152 10
rect 156 6 157 10
rect 148 3 157 6
rect 160 10 169 11
rect 160 6 161 10
rect 165 6 169 10
rect 160 3 169 6
rect 172 8 181 11
rect 172 4 176 8
rect 180 4 181 8
rect 172 3 181 4
rect 184 10 193 11
rect 184 6 185 10
rect 189 6 193 10
rect 184 3 193 6
rect 196 3 217 11
rect 220 10 229 11
rect 220 6 224 10
rect 228 6 229 10
rect 220 3 229 6
<< ndcontact >>
rect -133 -14 -129 -10
rect -94 -14 -90 -10
rect -85 -14 -81 -10
rect -46 -14 -42 -10
rect -37 -14 -33 -10
rect -22 -14 -18 -10
rect -10 -14 -6 -10
rect 29 -14 33 -10
rect 38 -14 42 -10
rect 77 -14 81 -10
rect 86 -14 90 -10
rect 101 -14 105 -10
rect 113 -14 117 -10
rect 152 -14 156 -10
rect 161 -14 165 -10
rect 200 -14 204 -10
rect 209 -14 213 -10
rect 224 -14 228 -10
<< pdcontact >>
rect -109 4 -105 8
rect -94 6 -90 10
rect -85 6 -81 10
rect -70 4 -66 8
rect -61 6 -57 10
rect -22 6 -18 10
rect 14 4 18 8
rect 29 6 33 10
rect 38 6 42 10
rect 53 4 57 8
rect 62 6 66 10
rect 101 6 105 10
rect 137 4 141 8
rect 152 6 156 10
rect 161 6 165 10
rect 176 4 180 8
rect 185 6 189 10
rect 224 6 228 10
<< psubstratepcontact >>
rect -130 -28 -126 -24
rect -122 -28 -118 -24
rect -114 -28 -110 -24
rect -106 -28 -102 -24
rect -98 -28 -94 -24
rect -90 -28 -86 -24
rect -82 -28 -78 -24
rect -74 -28 -70 -24
rect -66 -28 -62 -24
rect -58 -28 -54 -24
rect -50 -28 -46 -24
rect -42 -28 -38 -24
rect -34 -28 -30 -24
rect -26 -28 -22 -24
rect -18 -28 -14 -24
rect -7 -28 -3 -24
rect 1 -28 5 -24
rect 9 -28 13 -24
rect 17 -28 21 -24
rect 25 -28 29 -24
rect 33 -28 37 -24
rect 41 -28 45 -24
rect 49 -28 53 -24
rect 57 -28 61 -24
rect 65 -28 69 -24
rect 73 -28 77 -24
rect 81 -28 85 -24
rect 89 -28 93 -24
rect 97 -28 101 -24
rect 105 -28 109 -24
rect 116 -28 120 -24
rect 124 -28 128 -24
rect 132 -28 136 -24
rect 140 -28 144 -24
rect 148 -28 152 -24
rect 156 -28 160 -24
rect 164 -28 168 -24
rect 172 -28 176 -24
rect 180 -28 184 -24
rect 188 -28 192 -24
rect 196 -28 200 -24
rect 204 -28 208 -24
rect 212 -28 216 -24
rect 220 -28 224 -24
rect 228 -28 232 -24
<< nsubstratencontact >>
rect -131 20 -127 24
rect -123 20 -119 24
rect -115 20 -111 24
rect -107 20 -103 24
rect -99 20 -95 24
rect -91 20 -87 24
rect -83 20 -79 24
rect -75 20 -71 24
rect -67 20 -63 24
rect -59 20 -55 24
rect -51 20 -47 24
rect -43 20 -39 24
rect -35 20 -31 24
rect -27 20 -23 24
rect -19 20 -15 24
rect -8 20 -4 24
rect 0 20 4 24
rect 8 20 12 24
rect 16 20 20 24
rect 24 20 28 24
rect 32 20 36 24
rect 40 20 44 24
rect 48 20 52 24
rect 56 20 60 24
rect 64 20 68 24
rect 72 20 76 24
rect 80 20 84 24
rect 88 20 92 24
rect 96 20 100 24
rect 104 20 108 24
rect 115 20 119 24
rect 123 20 127 24
rect 131 20 135 24
rect 139 20 143 24
rect 147 20 151 24
rect 155 20 159 24
rect 163 20 167 24
rect 171 20 175 24
rect 179 20 183 24
rect 187 20 191 24
rect 195 20 199 24
rect 203 20 207 24
rect 211 20 215 24
rect 219 20 223 24
rect 227 20 231 24
<< polysilicon >>
rect -101 11 -98 13
rect -77 11 -74 13
rect -53 11 -50 12
rect -29 11 -26 13
rect 22 11 25 13
rect 46 11 49 13
rect 70 11 73 12
rect 94 11 97 13
rect 145 11 148 13
rect 169 11 172 13
rect 193 11 196 12
rect 217 11 220 13
rect -101 2 -98 3
rect -125 -9 -122 -7
rect -101 -9 -98 -2
rect -77 -9 -74 3
rect -53 2 -50 3
rect -29 1 -26 3
rect 22 2 25 3
rect -53 -9 -50 -7
rect -29 -9 -26 -7
rect -2 -9 1 -7
rect 22 -9 25 -2
rect 46 -9 49 3
rect 70 2 73 3
rect 94 1 97 3
rect 145 2 148 3
rect 70 -9 73 -7
rect 94 -9 97 -7
rect 121 -9 124 -7
rect 145 -9 148 -2
rect 169 -9 172 3
rect 193 2 196 3
rect 217 1 220 3
rect 193 -9 196 -7
rect 217 -9 220 -7
rect -125 -17 -122 -15
rect -101 -17 -98 -15
rect -77 -17 -74 -15
rect -53 -17 -50 -15
rect -29 -17 -26 -15
rect -2 -17 1 -15
rect 22 -17 25 -15
rect 46 -17 49 -15
rect 70 -17 73 -15
rect 94 -17 97 -15
rect 121 -17 124 -15
rect 145 -17 148 -15
rect 169 -17 172 -15
rect 193 -17 196 -15
rect 217 -17 220 -15
<< polycontact >>
rect -77 13 -73 17
rect -53 12 -49 16
rect -30 13 -26 17
rect 46 13 50 17
rect 70 12 74 16
rect 93 13 97 17
rect 169 13 173 17
rect 193 12 197 16
rect 216 13 220 17
rect -101 -2 -97 2
rect -125 -7 -121 -3
rect -54 -2 -50 2
rect 22 -2 26 2
rect -30 -7 -26 -3
rect -2 -7 2 -3
rect 69 -2 73 2
rect 145 -2 149 2
rect 93 -7 97 -3
rect 121 -7 125 -3
rect 192 -2 196 2
rect 216 -7 220 -3
rect -53 -21 -49 -17
rect 70 -21 74 -17
rect 193 -21 197 -17
<< metal1 >>
rect -134 20 -131 24
rect -127 20 -123 24
rect -119 20 -115 24
rect -111 20 -107 24
rect -103 20 -99 24
rect -95 20 -91 24
rect -87 20 -83 24
rect -79 20 -75 24
rect -71 20 -67 24
rect -63 20 -59 24
rect -55 20 -51 24
rect -47 20 -43 24
rect -39 20 -35 24
rect -31 20 -27 24
rect -23 20 -19 24
rect -15 20 -8 24
rect -4 20 0 24
rect 4 20 8 24
rect 12 20 16 24
rect 20 20 24 24
rect 28 20 32 24
rect 36 20 40 24
rect 44 20 48 24
rect 52 20 56 24
rect 60 20 64 24
rect 68 20 72 24
rect 76 20 80 24
rect 84 20 88 24
rect 92 20 96 24
rect 100 20 104 24
rect 108 20 115 24
rect 119 20 123 24
rect 127 20 131 24
rect 135 20 139 24
rect 143 20 147 24
rect 151 20 155 24
rect 159 20 163 24
rect 167 20 171 24
rect 175 20 179 24
rect 183 20 187 24
rect 191 20 195 24
rect 199 20 203 24
rect 207 20 211 24
rect 215 20 219 24
rect 223 20 227 24
rect 231 20 235 24
rect -134 13 -129 16
rect -132 7 -129 13
rect -93 10 -90 20
rect -132 4 -109 7
rect -85 10 -82 20
rect -73 13 -72 17
rect -60 10 -57 20
rect -49 12 -39 15
rect -31 13 -30 17
rect -26 13 -6 16
rect -132 -10 -129 4
rect -69 1 -66 4
rect -97 -2 -66 1
rect -55 -2 -54 2
rect -125 -3 -121 -2
rect -69 -10 -66 -2
rect -42 -3 -39 12
rect -42 -6 -30 -3
rect -21 -10 -18 6
rect -9 7 -6 13
rect 30 10 33 20
rect -9 4 14 7
rect 38 10 41 20
rect 50 13 51 17
rect 63 10 66 20
rect 74 12 84 15
rect 92 13 93 17
rect 97 13 117 16
rect -9 -10 -6 4
rect 54 1 57 4
rect 26 -2 57 1
rect 68 -2 69 2
rect -2 -3 2 -2
rect 54 -10 57 -2
rect 81 -3 84 12
rect 81 -6 93 -3
rect 102 -10 105 6
rect 114 7 117 13
rect 153 10 156 20
rect 114 4 137 7
rect 161 10 164 20
rect 173 13 174 17
rect 186 10 189 20
rect 197 12 207 15
rect 215 13 216 17
rect 220 13 235 16
rect 114 -10 117 4
rect 177 1 180 4
rect 149 -2 180 1
rect 191 -2 192 2
rect 121 -3 125 -2
rect 177 -10 180 -2
rect 204 -3 207 12
rect 204 -6 216 -3
rect 225 -10 228 6
rect -93 -24 -90 -14
rect -69 -13 -46 -10
rect -85 -24 -82 -14
rect -49 -21 -48 -17
rect -37 -24 -34 -14
rect 30 -24 33 -14
rect 54 -13 77 -10
rect 38 -24 41 -14
rect 74 -21 75 -17
rect 86 -24 89 -14
rect 153 -24 156 -14
rect 177 -13 200 -10
rect 161 -24 164 -14
rect 197 -21 198 -17
rect 209 -24 212 -14
rect -134 -28 -130 -24
rect -126 -28 -122 -24
rect -118 -28 -114 -24
rect -110 -28 -106 -24
rect -102 -28 -98 -24
rect -94 -28 -90 -24
rect -86 -28 -82 -24
rect -78 -28 -74 -24
rect -70 -28 -66 -24
rect -62 -28 -58 -24
rect -54 -28 -50 -24
rect -46 -28 -42 -24
rect -38 -28 -34 -24
rect -30 -28 -26 -24
rect -22 -28 -18 -24
rect -14 -28 -7 -24
rect -3 -28 1 -24
rect 5 -28 9 -24
rect 13 -28 17 -24
rect 21 -28 25 -24
rect 29 -28 33 -24
rect 37 -28 41 -24
rect 45 -28 49 -24
rect 53 -28 57 -24
rect 61 -28 65 -24
rect 69 -28 73 -24
rect 77 -28 81 -24
rect 85 -28 89 -24
rect 93 -28 97 -24
rect 101 -28 105 -24
rect 109 -28 116 -24
rect 120 -28 124 -24
rect 128 -28 132 -24
rect 136 -28 140 -24
rect 144 -28 148 -24
rect 152 -28 156 -24
rect 160 -28 164 -24
rect 168 -28 172 -24
rect 176 -28 180 -24
rect 184 -28 188 -24
rect 192 -28 196 -24
rect 200 -28 204 -24
rect 208 -28 212 -24
rect 216 -28 220 -24
rect 224 -28 228 -24
rect 232 -28 235 -24
<< m2contact >>
rect -77 13 -73 17
rect -30 13 -26 17
rect -54 -2 -50 2
rect -125 -7 -121 -3
rect 46 13 50 17
rect 93 13 97 17
rect 69 -2 73 2
rect -2 -7 2 -3
rect 169 13 173 17
rect 216 13 220 17
rect 192 -2 196 2
rect 121 -7 125 -3
rect -133 -14 -129 -10
rect -22 -14 -18 -10
rect -10 -14 -6 -10
rect -53 -21 -49 -17
rect 101 -14 105 -10
rect 113 -14 117 -10
rect 70 -21 74 -17
rect 224 -14 228 -10
rect 193 -21 197 -17
<< metal2 >>
rect -125 13 -77 16
rect -73 13 -30 16
rect -2 13 46 16
rect 50 13 93 16
rect 121 13 169 16
rect 173 13 216 16
rect -125 -3 -122 13
rect -53 -10 -50 -2
rect -2 -3 1 13
rect 70 -10 73 -2
rect 121 -3 124 13
rect 193 -10 196 -2
rect -129 -13 -50 -10
rect -6 -13 73 -10
rect 117 -13 196 -10
rect -22 -18 -19 -14
rect -49 -21 -19 -18
rect 101 -18 104 -14
rect 74 -21 104 -18
rect 224 -18 227 -14
rect 197 -21 227 -18
<< labels >>
rlabel metal1 -134 13 -134 16 3 out
rlabel metal1 -132 22 -132 22 4 vdd!
rlabel metal1 -132 -26 -132 -26 2 gnd!
rlabel metal1 235 13 235 16 7 in
<< end >>
