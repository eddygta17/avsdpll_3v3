magic
tech scmos
timestamp 1599387223
<< nwell >>
rect -11 -3 112 27
<< ntransistor >>
rect -2 -15 1 -9
rect 22 -15 25 -9
rect 46 -15 49 -9
rect 70 -15 73 -9
rect 94 -15 97 -9
<< ptransistor >>
rect 22 3 25 11
rect 46 3 49 11
rect 70 3 73 11
rect 94 3 97 11
<< ndiffusion >>
rect -11 -10 -2 -9
rect -11 -14 -10 -10
rect -6 -14 -2 -10
rect -11 -15 -2 -14
rect 1 -15 22 -9
rect 25 -10 34 -9
rect 25 -14 29 -10
rect 33 -14 34 -10
rect 25 -15 34 -14
rect 37 -10 46 -9
rect 37 -14 38 -10
rect 42 -14 46 -10
rect 37 -15 46 -14
rect 49 -15 70 -9
rect 73 -10 82 -9
rect 73 -14 77 -10
rect 81 -14 82 -10
rect 73 -15 82 -14
rect 85 -10 94 -9
rect 85 -14 86 -10
rect 90 -14 94 -10
rect 85 -15 94 -14
rect 97 -10 106 -9
rect 97 -14 101 -10
rect 105 -14 106 -10
rect 97 -15 106 -14
<< pdiffusion >>
rect 13 8 22 11
rect 13 4 14 8
rect 18 4 22 8
rect 13 3 22 4
rect 25 10 34 11
rect 25 6 29 10
rect 33 6 34 10
rect 25 3 34 6
rect 37 10 46 11
rect 37 6 38 10
rect 42 6 46 10
rect 37 3 46 6
rect 49 8 58 11
rect 49 4 53 8
rect 57 4 58 8
rect 49 3 58 4
rect 61 10 70 11
rect 61 6 62 10
rect 66 6 70 10
rect 61 3 70 6
rect 73 3 94 11
rect 97 10 106 11
rect 97 6 101 10
rect 105 6 106 10
rect 97 3 106 6
<< ndcontact >>
rect -10 -14 -6 -10
rect 29 -14 33 -10
rect 38 -14 42 -10
rect 77 -14 81 -10
rect 86 -14 90 -10
rect 101 -14 105 -10
<< pdcontact >>
rect 14 4 18 8
rect 29 6 33 10
rect 38 6 42 10
rect 53 4 57 8
rect 62 6 66 10
rect 101 6 105 10
<< psubstratepcontact >>
rect -7 -28 -3 -24
rect 1 -28 5 -24
rect 9 -28 13 -24
rect 17 -28 21 -24
rect 25 -28 29 -24
rect 33 -28 37 -24
rect 41 -28 45 -24
rect 49 -28 53 -24
rect 57 -28 61 -24
rect 65 -28 69 -24
rect 73 -28 77 -24
rect 81 -28 85 -24
rect 89 -28 93 -24
rect 97 -28 101 -24
rect 105 -28 109 -24
<< nsubstratencontact >>
rect -8 20 -4 24
rect 0 20 4 24
rect 8 20 12 24
rect 16 20 20 24
rect 24 20 28 24
rect 32 20 36 24
rect 40 20 44 24
rect 48 20 52 24
rect 56 20 60 24
rect 64 20 68 24
rect 72 20 76 24
rect 80 20 84 24
rect 88 20 92 24
rect 96 20 100 24
rect 104 20 108 24
<< polysilicon >>
rect 22 11 25 13
rect 46 11 49 13
rect 70 11 73 12
rect 94 11 97 13
rect 22 2 25 3
rect -2 -9 1 -7
rect 22 -9 25 -2
rect 46 -9 49 3
rect 70 2 73 3
rect 94 1 97 3
rect 70 -9 73 -7
rect 94 -9 97 -7
rect -2 -17 1 -15
rect 22 -17 25 -15
rect 46 -17 49 -15
rect 70 -17 73 -15
rect 94 -17 97 -15
<< polycontact >>
rect 46 13 50 17
rect 70 12 74 16
rect 93 13 97 17
rect 22 -2 26 2
rect -2 -7 2 -3
rect 69 -2 73 2
rect 93 -7 97 -3
rect 70 -21 74 -17
<< metal1 >>
rect -11 20 -8 24
rect -4 20 0 24
rect 4 20 8 24
rect 12 20 16 24
rect 20 20 24 24
rect 28 20 32 24
rect 36 20 40 24
rect 44 20 48 24
rect 52 20 56 24
rect 60 20 64 24
rect 68 20 72 24
rect 76 20 80 24
rect 84 20 88 24
rect 92 20 96 24
rect 100 20 104 24
rect 108 20 112 24
rect -11 13 -6 16
rect -9 7 -6 13
rect 30 10 33 20
rect -9 4 14 7
rect 38 10 41 20
rect 50 13 51 17
rect 63 10 66 20
rect 74 12 84 15
rect 92 13 93 17
rect 97 13 112 16
rect -9 -10 -6 4
rect 54 1 57 4
rect 26 -2 57 1
rect 68 -2 69 2
rect -2 -3 2 -2
rect 54 -10 57 -2
rect 81 -3 84 12
rect 81 -6 93 -3
rect 102 -10 105 6
rect 30 -24 33 -14
rect 54 -13 77 -10
rect 38 -24 41 -14
rect 74 -21 75 -17
rect 86 -24 89 -14
rect -11 -28 -7 -24
rect -3 -28 1 -24
rect 5 -28 9 -24
rect 13 -28 17 -24
rect 21 -28 25 -24
rect 29 -28 33 -24
rect 37 -28 41 -24
rect 45 -28 49 -24
rect 53 -28 57 -24
rect 61 -28 65 -24
rect 69 -28 73 -24
rect 77 -28 81 -24
rect 85 -28 89 -24
rect 93 -28 97 -24
rect 101 -28 105 -24
rect 109 -28 112 -24
<< m2contact >>
rect 46 13 50 17
rect 93 13 97 17
rect 69 -2 73 2
rect -2 -7 2 -3
rect -10 -14 -6 -10
rect 101 -14 105 -10
rect 70 -21 74 -17
<< metal2 >>
rect -2 13 46 16
rect 50 13 93 16
rect -2 -3 1 13
rect 70 -10 73 -2
rect -6 -13 73 -10
rect 101 -18 104 -14
rect 74 -21 104 -18
<< labels >>
rlabel metal1 -9 22 -9 22 4 vdd!
rlabel metal1 -8 -26 -8 -26 2 gnd!
rlabel metal1 -11 13 -11 16 3 out
rlabel metal1 112 13 112 16 7 in
<< end >>
