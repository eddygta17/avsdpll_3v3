magic
tech scmos
timestamp 1599410049
<< nwell >>
rect 27 150 913 207
rect 27 -11 876 46
<< ntransistor >>
rect 48 108 50 128
rect 53 108 55 128
rect 69 108 71 128
rect 74 108 76 128
rect 104 108 106 128
rect 109 108 111 128
rect 125 108 127 128
rect 130 108 132 128
rect 160 108 162 128
rect 165 108 167 128
rect 181 108 183 128
rect 186 108 188 128
rect 216 108 218 128
rect 221 108 223 128
rect 237 108 239 128
rect 242 108 244 128
rect 272 108 274 128
rect 277 108 279 128
rect 293 108 295 128
rect 298 108 300 128
rect 328 108 330 128
rect 333 108 335 128
rect 349 108 351 128
rect 354 108 356 128
rect 384 108 386 128
rect 389 108 391 128
rect 405 108 407 128
rect 410 108 412 128
rect 440 108 442 128
rect 445 108 447 128
rect 461 108 463 128
rect 466 108 468 128
rect 496 108 498 128
rect 501 108 503 128
rect 517 108 519 128
rect 522 108 524 128
rect 552 108 554 128
rect 557 108 559 128
rect 573 108 575 128
rect 578 108 580 128
rect 608 108 610 128
rect 613 108 615 128
rect 629 108 631 128
rect 634 108 636 128
rect 664 108 666 128
rect 669 108 671 128
rect 685 108 687 128
rect 690 108 692 128
rect 720 108 722 128
rect 725 108 727 128
rect 741 108 743 128
rect 746 108 748 128
rect 776 108 778 128
rect 781 108 783 128
rect 797 108 799 128
rect 802 108 804 128
rect 832 108 834 128
rect 837 108 839 128
rect 853 108 855 128
rect 858 108 860 128
rect 892 108 894 128
rect 900 108 902 128
rect 48 68 50 88
rect 53 68 55 88
rect 69 68 71 88
rect 74 68 76 88
rect 104 68 106 88
rect 109 68 111 88
rect 125 68 127 88
rect 130 68 132 88
rect 160 68 162 88
rect 165 68 167 88
rect 181 68 183 88
rect 186 68 188 88
rect 216 68 218 88
rect 221 68 223 88
rect 237 68 239 88
rect 242 68 244 88
rect 272 68 274 88
rect 277 68 279 88
rect 293 68 295 88
rect 298 68 300 88
rect 328 68 330 88
rect 333 68 335 88
rect 349 68 351 88
rect 354 68 356 88
rect 384 68 386 88
rect 389 68 391 88
rect 405 68 407 88
rect 410 68 412 88
rect 440 68 442 88
rect 445 68 447 88
rect 461 68 463 88
rect 466 68 468 88
rect 496 68 498 88
rect 501 68 503 88
rect 517 68 519 88
rect 522 68 524 88
rect 552 68 554 88
rect 557 68 559 88
rect 573 68 575 88
rect 578 68 580 88
rect 608 68 610 88
rect 613 68 615 88
rect 629 68 631 88
rect 634 68 636 88
rect 664 68 666 88
rect 669 68 671 88
rect 685 68 687 88
rect 690 68 692 88
rect 720 68 722 88
rect 725 68 727 88
rect 741 68 743 88
rect 746 68 748 88
rect 776 68 778 88
rect 781 68 783 88
rect 797 68 799 88
rect 802 68 804 88
rect 832 68 834 88
rect 837 68 839 88
rect 853 68 855 88
rect 858 68 860 88
<< ptransistor >>
rect 53 156 55 196
rect 74 156 76 196
rect 109 156 111 196
rect 130 156 132 196
rect 165 156 167 196
rect 186 156 188 196
rect 221 156 223 196
rect 242 156 244 196
rect 277 156 279 196
rect 298 156 300 196
rect 333 156 335 196
rect 354 156 356 196
rect 389 156 391 196
rect 410 156 412 196
rect 445 156 447 196
rect 466 156 468 196
rect 501 156 503 196
rect 522 156 524 196
rect 557 156 559 196
rect 578 156 580 196
rect 613 156 615 196
rect 634 156 636 196
rect 669 156 671 196
rect 690 156 692 196
rect 725 156 727 196
rect 746 156 748 196
rect 781 156 783 196
rect 802 156 804 196
rect 837 156 839 196
rect 858 156 860 196
rect 892 156 894 196
rect 900 156 902 196
rect 53 0 55 40
rect 74 0 76 40
rect 109 0 111 40
rect 130 0 132 40
rect 165 0 167 40
rect 186 0 188 40
rect 221 0 223 40
rect 242 0 244 40
rect 277 0 279 40
rect 298 0 300 40
rect 333 0 335 40
rect 354 0 356 40
rect 389 0 391 40
rect 410 0 412 40
rect 445 0 447 40
rect 466 0 468 40
rect 501 0 503 40
rect 522 0 524 40
rect 557 0 559 40
rect 578 0 580 40
rect 613 0 615 40
rect 634 0 636 40
rect 669 0 671 40
rect 690 0 692 40
rect 725 0 727 40
rect 746 0 748 40
rect 781 0 783 40
rect 802 0 804 40
rect 837 0 839 40
rect 858 0 860 40
<< ndiffusion >>
rect 47 108 48 128
rect 50 108 53 128
rect 55 108 56 128
rect 68 108 69 128
rect 71 108 74 128
rect 76 108 77 128
rect 103 108 104 128
rect 106 108 109 128
rect 111 108 112 128
rect 124 108 125 128
rect 127 108 130 128
rect 132 108 133 128
rect 159 108 160 128
rect 162 108 165 128
rect 167 108 168 128
rect 180 108 181 128
rect 183 108 186 128
rect 188 108 189 128
rect 215 108 216 128
rect 218 108 221 128
rect 223 108 224 128
rect 236 108 237 128
rect 239 108 242 128
rect 244 108 245 128
rect 271 108 272 128
rect 274 108 277 128
rect 279 108 280 128
rect 292 108 293 128
rect 295 108 298 128
rect 300 108 301 128
rect 327 108 328 128
rect 330 108 333 128
rect 335 108 336 128
rect 348 108 349 128
rect 351 108 354 128
rect 356 108 357 128
rect 383 108 384 128
rect 386 108 389 128
rect 391 108 392 128
rect 404 108 405 128
rect 407 108 410 128
rect 412 108 413 128
rect 439 108 440 128
rect 442 108 445 128
rect 447 108 448 128
rect 460 108 461 128
rect 463 108 466 128
rect 468 108 469 128
rect 495 108 496 128
rect 498 108 501 128
rect 503 108 504 128
rect 516 108 517 128
rect 519 108 522 128
rect 524 108 525 128
rect 551 108 552 128
rect 554 108 557 128
rect 559 108 560 128
rect 572 108 573 128
rect 575 108 578 128
rect 580 108 581 128
rect 607 108 608 128
rect 610 108 613 128
rect 615 108 616 128
rect 628 108 629 128
rect 631 108 634 128
rect 636 108 637 128
rect 663 108 664 128
rect 666 108 669 128
rect 671 108 672 128
rect 684 108 685 128
rect 687 108 690 128
rect 692 108 693 128
rect 719 108 720 128
rect 722 108 725 128
rect 727 108 728 128
rect 740 108 741 128
rect 743 108 746 128
rect 748 108 749 128
rect 775 108 776 128
rect 778 108 781 128
rect 783 108 784 128
rect 796 108 797 128
rect 799 108 802 128
rect 804 108 805 128
rect 831 108 832 128
rect 834 108 837 128
rect 839 108 840 128
rect 852 108 853 128
rect 855 108 858 128
rect 860 108 861 128
rect 891 108 892 128
rect 894 108 895 128
rect 899 108 900 128
rect 902 108 903 128
rect 47 68 48 88
rect 50 68 53 88
rect 55 68 56 88
rect 68 68 69 88
rect 71 68 74 88
rect 76 68 77 88
rect 103 68 104 88
rect 106 68 109 88
rect 111 68 112 88
rect 124 68 125 88
rect 127 68 130 88
rect 132 68 133 88
rect 159 68 160 88
rect 162 68 165 88
rect 167 68 168 88
rect 180 68 181 88
rect 183 68 186 88
rect 188 68 189 88
rect 215 68 216 88
rect 218 68 221 88
rect 223 68 224 88
rect 236 68 237 88
rect 239 68 242 88
rect 244 68 245 88
rect 271 68 272 88
rect 274 68 277 88
rect 279 68 280 88
rect 292 68 293 88
rect 295 68 298 88
rect 300 68 301 88
rect 327 68 328 88
rect 330 68 333 88
rect 335 68 336 88
rect 348 68 349 88
rect 351 68 354 88
rect 356 68 357 88
rect 383 68 384 88
rect 386 68 389 88
rect 391 68 392 88
rect 404 68 405 88
rect 407 68 410 88
rect 412 68 413 88
rect 439 68 440 88
rect 442 68 445 88
rect 447 68 448 88
rect 460 68 461 88
rect 463 68 466 88
rect 468 68 469 88
rect 495 68 496 88
rect 498 68 501 88
rect 503 68 504 88
rect 516 68 517 88
rect 519 68 522 88
rect 524 68 525 88
rect 551 68 552 88
rect 554 68 557 88
rect 559 68 560 88
rect 572 68 573 88
rect 575 68 578 88
rect 580 68 581 88
rect 607 68 608 88
rect 610 68 613 88
rect 615 68 616 88
rect 628 68 629 88
rect 631 68 634 88
rect 636 68 637 88
rect 663 68 664 88
rect 666 68 669 88
rect 671 68 672 88
rect 684 68 685 88
rect 687 68 690 88
rect 692 68 693 88
rect 719 68 720 88
rect 722 68 725 88
rect 727 68 728 88
rect 740 68 741 88
rect 743 68 746 88
rect 748 68 749 88
rect 775 68 776 88
rect 778 68 781 88
rect 783 68 784 88
rect 796 68 797 88
rect 799 68 802 88
rect 804 68 805 88
rect 831 68 832 88
rect 834 68 837 88
rect 839 68 840 88
rect 852 68 853 88
rect 855 68 858 88
rect 860 68 861 88
<< pdiffusion >>
rect 52 156 53 196
rect 55 156 56 196
rect 73 156 74 196
rect 76 156 77 196
rect 108 156 109 196
rect 111 156 112 196
rect 129 156 130 196
rect 132 156 133 196
rect 164 156 165 196
rect 167 156 168 196
rect 185 156 186 196
rect 188 156 189 196
rect 220 156 221 196
rect 223 156 224 196
rect 241 156 242 196
rect 244 156 245 196
rect 276 156 277 196
rect 279 156 280 196
rect 297 156 298 196
rect 300 156 301 196
rect 332 156 333 196
rect 335 156 336 196
rect 353 156 354 196
rect 356 156 357 196
rect 388 156 389 196
rect 391 156 392 196
rect 409 156 410 196
rect 412 156 413 196
rect 444 156 445 196
rect 447 156 448 196
rect 465 156 466 196
rect 468 156 469 196
rect 500 156 501 196
rect 503 156 504 196
rect 521 156 522 196
rect 524 156 525 196
rect 556 156 557 196
rect 559 156 560 196
rect 577 156 578 196
rect 580 156 581 196
rect 612 156 613 196
rect 615 156 616 196
rect 633 156 634 196
rect 636 156 637 196
rect 668 156 669 196
rect 671 156 672 196
rect 689 156 690 196
rect 692 156 693 196
rect 724 156 725 196
rect 727 156 728 196
rect 745 156 746 196
rect 748 156 749 196
rect 780 156 781 196
rect 783 156 784 196
rect 801 156 802 196
rect 804 156 805 196
rect 836 156 837 196
rect 839 156 840 196
rect 857 156 858 196
rect 860 156 861 196
rect 891 156 892 196
rect 894 156 895 196
rect 899 156 900 196
rect 902 156 903 196
rect 52 0 53 40
rect 55 0 56 40
rect 73 0 74 40
rect 76 0 77 40
rect 108 0 109 40
rect 111 0 112 40
rect 129 0 130 40
rect 132 0 133 40
rect 164 0 165 40
rect 167 0 168 40
rect 185 0 186 40
rect 188 0 189 40
rect 220 0 221 40
rect 223 0 224 40
rect 241 0 242 40
rect 244 0 245 40
rect 276 0 277 40
rect 279 0 280 40
rect 297 0 298 40
rect 300 0 301 40
rect 332 0 333 40
rect 335 0 336 40
rect 353 0 354 40
rect 356 0 357 40
rect 388 0 389 40
rect 391 0 392 40
rect 409 0 410 40
rect 412 0 413 40
rect 444 0 445 40
rect 447 0 448 40
rect 465 0 466 40
rect 468 0 469 40
rect 500 0 501 40
rect 503 0 504 40
rect 521 0 522 40
rect 524 0 525 40
rect 556 0 557 40
rect 559 0 560 40
rect 577 0 578 40
rect 580 0 581 40
rect 612 0 613 40
rect 615 0 616 40
rect 633 0 634 40
rect 636 0 637 40
rect 668 0 669 40
rect 671 0 672 40
rect 689 0 690 40
rect 692 0 693 40
rect 724 0 725 40
rect 727 0 728 40
rect 745 0 746 40
rect 748 0 749 40
rect 780 0 781 40
rect 783 0 784 40
rect 801 0 802 40
rect 804 0 805 40
rect 836 0 837 40
rect 839 0 840 40
rect 857 0 858 40
rect 860 0 861 40
<< ndcontact >>
rect 43 108 47 128
rect 56 108 60 128
rect 64 108 68 128
rect 77 108 81 128
rect 99 108 103 128
rect 112 108 116 128
rect 120 108 124 128
rect 133 108 137 128
rect 155 108 159 128
rect 168 108 172 128
rect 176 108 180 128
rect 189 108 193 128
rect 211 108 215 128
rect 224 108 228 128
rect 232 108 236 128
rect 245 108 249 128
rect 267 108 271 128
rect 280 108 284 128
rect 288 108 292 128
rect 301 108 305 128
rect 323 108 327 128
rect 336 108 340 128
rect 344 108 348 128
rect 357 108 361 128
rect 379 108 383 128
rect 392 108 396 128
rect 400 108 404 128
rect 413 108 417 128
rect 435 108 439 128
rect 448 108 452 128
rect 456 108 460 128
rect 469 108 473 128
rect 491 108 495 128
rect 504 108 508 128
rect 512 108 516 128
rect 525 108 529 128
rect 547 108 551 128
rect 560 108 564 128
rect 568 108 572 128
rect 581 108 585 128
rect 603 108 607 128
rect 616 108 620 128
rect 624 108 628 128
rect 637 108 641 128
rect 659 108 663 128
rect 672 108 676 128
rect 680 108 684 128
rect 693 108 697 128
rect 715 108 719 128
rect 728 108 732 128
rect 736 108 740 128
rect 749 108 753 128
rect 771 108 775 128
rect 784 108 788 128
rect 792 108 796 128
rect 805 108 809 128
rect 827 108 831 128
rect 840 108 844 128
rect 848 108 852 128
rect 861 108 865 128
rect 887 108 891 128
rect 895 108 899 128
rect 903 108 907 128
rect 43 68 47 88
rect 56 68 60 88
rect 64 68 68 88
rect 77 68 81 88
rect 99 68 103 88
rect 112 68 116 88
rect 120 68 124 88
rect 133 68 137 88
rect 155 68 159 88
rect 168 68 172 88
rect 176 68 180 88
rect 189 68 193 88
rect 211 68 215 88
rect 224 68 228 88
rect 232 68 236 88
rect 245 68 249 88
rect 267 68 271 88
rect 280 68 284 88
rect 288 68 292 88
rect 301 68 305 88
rect 323 68 327 88
rect 336 68 340 88
rect 344 68 348 88
rect 357 68 361 88
rect 379 68 383 88
rect 392 68 396 88
rect 400 68 404 88
rect 413 68 417 88
rect 435 68 439 88
rect 448 68 452 88
rect 456 68 460 88
rect 469 68 473 88
rect 491 68 495 88
rect 504 68 508 88
rect 512 68 516 88
rect 525 68 529 88
rect 547 68 551 88
rect 560 68 564 88
rect 568 68 572 88
rect 581 68 585 88
rect 603 68 607 88
rect 616 68 620 88
rect 624 68 628 88
rect 637 68 641 88
rect 659 68 663 88
rect 672 68 676 88
rect 680 68 684 88
rect 693 68 697 88
rect 715 68 719 88
rect 728 68 732 88
rect 736 68 740 88
rect 749 68 753 88
rect 771 68 775 88
rect 784 68 788 88
rect 792 68 796 88
rect 805 68 809 88
rect 827 68 831 88
rect 840 68 844 88
rect 848 68 852 88
rect 861 68 865 88
<< pdcontact >>
rect 48 156 52 196
rect 56 156 60 196
rect 69 156 73 196
rect 77 156 81 196
rect 104 156 108 196
rect 112 156 116 196
rect 125 156 129 196
rect 133 156 137 196
rect 160 156 164 196
rect 168 156 172 196
rect 181 156 185 196
rect 189 156 193 196
rect 216 156 220 196
rect 224 156 228 196
rect 237 156 241 196
rect 245 156 249 196
rect 272 156 276 196
rect 280 156 284 196
rect 293 156 297 196
rect 301 156 305 196
rect 328 156 332 196
rect 336 156 340 196
rect 349 156 353 196
rect 357 156 361 196
rect 384 156 388 196
rect 392 156 396 196
rect 405 156 409 196
rect 413 156 417 196
rect 440 156 444 196
rect 448 156 452 196
rect 461 156 465 196
rect 469 156 473 196
rect 496 156 500 196
rect 504 156 508 196
rect 517 156 521 196
rect 525 156 529 196
rect 552 156 556 196
rect 560 156 564 196
rect 573 156 577 196
rect 581 156 585 196
rect 608 156 612 196
rect 616 156 620 196
rect 629 156 633 196
rect 637 156 641 196
rect 664 156 668 196
rect 672 156 676 196
rect 685 156 689 196
rect 693 156 697 196
rect 720 156 724 196
rect 728 156 732 196
rect 741 156 745 196
rect 749 156 753 196
rect 776 156 780 196
rect 784 156 788 196
rect 797 156 801 196
rect 805 156 809 196
rect 832 156 836 196
rect 840 156 844 196
rect 853 156 857 196
rect 861 156 865 196
rect 887 156 891 196
rect 895 156 899 196
rect 903 156 907 196
rect 48 0 52 40
rect 56 0 60 40
rect 69 0 73 40
rect 77 0 81 40
rect 104 0 108 40
rect 112 0 116 40
rect 125 0 129 40
rect 133 0 137 40
rect 160 0 164 40
rect 168 0 172 40
rect 181 0 185 40
rect 189 0 193 40
rect 216 0 220 40
rect 224 0 228 40
rect 237 0 241 40
rect 245 0 249 40
rect 272 0 276 40
rect 280 0 284 40
rect 293 0 297 40
rect 301 0 305 40
rect 328 0 332 40
rect 336 0 340 40
rect 349 0 353 40
rect 357 0 361 40
rect 384 0 388 40
rect 392 0 396 40
rect 405 0 409 40
rect 413 0 417 40
rect 440 0 444 40
rect 448 0 452 40
rect 461 0 465 40
rect 469 0 473 40
rect 496 0 500 40
rect 504 0 508 40
rect 517 0 521 40
rect 525 0 529 40
rect 552 0 556 40
rect 560 0 564 40
rect 573 0 577 40
rect 581 0 585 40
rect 608 0 612 40
rect 616 0 620 40
rect 629 0 633 40
rect 637 0 641 40
rect 664 0 668 40
rect 672 0 676 40
rect 685 0 689 40
rect 693 0 697 40
rect 720 0 724 40
rect 728 0 732 40
rect 741 0 745 40
rect 749 0 753 40
rect 776 0 780 40
rect 784 0 788 40
rect 797 0 801 40
rect 805 0 809 40
rect 832 0 836 40
rect 840 0 844 40
rect 853 0 857 40
rect 861 0 865 40
<< psubstratepcontact >>
rect 51 100 55 104
rect 60 100 64 104
rect 72 100 76 104
rect 81 100 85 104
rect 98 100 102 104
rect 107 100 111 104
rect 116 100 120 104
rect 128 100 132 104
rect 137 100 141 104
rect 154 100 158 104
rect 163 100 167 104
rect 172 100 176 104
rect 184 100 188 104
rect 193 100 197 104
rect 210 100 214 104
rect 219 100 223 104
rect 228 100 232 104
rect 240 100 244 104
rect 249 100 253 104
rect 266 100 270 104
rect 275 100 279 104
rect 284 100 288 104
rect 296 100 300 104
rect 305 100 309 104
rect 322 100 326 104
rect 331 100 335 104
rect 340 100 344 104
rect 352 100 356 104
rect 361 100 365 104
rect 378 100 382 104
rect 387 100 391 104
rect 396 100 400 104
rect 408 100 412 104
rect 417 100 421 104
rect 434 100 438 104
rect 443 100 447 104
rect 452 100 456 104
rect 464 100 468 104
rect 473 100 477 104
rect 490 100 494 104
rect 499 100 503 104
rect 508 100 512 104
rect 520 100 524 104
rect 529 100 533 104
rect 546 100 550 104
rect 555 100 559 104
rect 564 100 568 104
rect 576 100 580 104
rect 585 100 589 104
rect 602 100 606 104
rect 611 100 615 104
rect 620 100 624 104
rect 632 100 636 104
rect 641 100 645 104
rect 658 100 662 104
rect 667 100 671 104
rect 676 100 680 104
rect 688 100 692 104
rect 697 100 701 104
rect 714 100 718 104
rect 723 100 727 104
rect 732 100 736 104
rect 744 100 748 104
rect 753 100 757 104
rect 770 100 774 104
rect 779 100 783 104
rect 788 100 792 104
rect 800 100 804 104
rect 809 100 813 104
rect 826 100 830 104
rect 835 100 839 104
rect 844 100 848 104
rect 856 100 860 104
rect 868 100 872 104
rect 883 100 887 104
rect 899 100 903 104
rect 51 92 55 96
rect 60 92 64 96
rect 72 92 76 96
rect 81 92 85 96
rect 98 92 102 96
rect 107 92 111 96
rect 116 92 120 96
rect 128 92 132 96
rect 137 92 141 96
rect 154 92 158 96
rect 163 92 167 96
rect 172 92 176 96
rect 184 92 188 96
rect 193 92 197 96
rect 210 92 214 96
rect 219 92 223 96
rect 228 92 232 96
rect 240 92 244 96
rect 249 92 253 96
rect 266 92 270 96
rect 275 92 279 96
rect 284 92 288 96
rect 296 92 300 96
rect 305 92 309 96
rect 322 92 326 96
rect 331 92 335 96
rect 340 92 344 96
rect 352 92 356 96
rect 361 92 365 96
rect 378 92 382 96
rect 387 92 391 96
rect 396 92 400 96
rect 408 92 412 96
rect 417 92 421 96
rect 434 92 438 96
rect 443 92 447 96
rect 452 92 456 96
rect 464 92 468 96
rect 473 92 477 96
rect 490 92 494 96
rect 499 92 503 96
rect 508 92 512 96
rect 520 92 524 96
rect 529 92 533 96
rect 546 92 550 96
rect 555 92 559 96
rect 564 92 568 96
rect 576 92 580 96
rect 585 92 589 96
rect 602 92 606 96
rect 611 92 615 96
rect 620 92 624 96
rect 632 92 636 96
rect 641 92 645 96
rect 658 92 662 96
rect 667 92 671 96
rect 676 92 680 96
rect 688 92 692 96
rect 697 92 701 96
rect 714 92 718 96
rect 723 92 727 96
rect 732 92 736 96
rect 744 92 748 96
rect 753 92 757 96
rect 770 92 774 96
rect 779 92 783 96
rect 788 92 792 96
rect 800 92 804 96
rect 809 92 813 96
rect 826 92 830 96
rect 835 92 839 96
rect 844 92 848 96
rect 856 92 860 96
rect 868 92 872 96
rect 883 92 887 96
rect 899 92 903 96
<< nsubstratencontact >>
rect 42 200 46 204
rect 51 200 55 204
rect 60 200 64 204
rect 72 200 76 204
rect 81 200 85 204
rect 98 200 102 204
rect 107 200 111 204
rect 116 200 120 204
rect 128 200 132 204
rect 137 200 141 204
rect 154 200 158 204
rect 163 200 167 204
rect 172 200 176 204
rect 184 200 188 204
rect 193 200 197 204
rect 210 200 214 204
rect 219 200 223 204
rect 228 200 232 204
rect 240 200 244 204
rect 249 200 253 204
rect 266 200 270 204
rect 275 200 279 204
rect 284 200 288 204
rect 296 200 300 204
rect 305 200 309 204
rect 322 200 326 204
rect 331 200 335 204
rect 340 200 344 204
rect 352 200 356 204
rect 361 200 365 204
rect 378 200 382 204
rect 387 200 391 204
rect 396 200 400 204
rect 408 200 412 204
rect 417 200 421 204
rect 434 200 438 204
rect 443 200 447 204
rect 452 200 456 204
rect 464 200 468 204
rect 473 200 477 204
rect 490 200 494 204
rect 499 200 503 204
rect 508 200 512 204
rect 520 200 524 204
rect 529 200 533 204
rect 546 200 550 204
rect 555 200 559 204
rect 564 200 568 204
rect 576 200 580 204
rect 585 200 589 204
rect 602 200 606 204
rect 611 200 615 204
rect 620 200 624 204
rect 632 200 636 204
rect 641 200 645 204
rect 658 200 662 204
rect 667 200 671 204
rect 676 200 680 204
rect 688 200 692 204
rect 697 200 701 204
rect 714 200 718 204
rect 723 200 727 204
rect 732 200 736 204
rect 744 200 748 204
rect 753 200 757 204
rect 770 200 774 204
rect 779 200 783 204
rect 788 200 792 204
rect 800 200 804 204
rect 809 200 813 204
rect 826 200 830 204
rect 835 200 839 204
rect 844 200 848 204
rect 856 200 860 204
rect 865 200 869 204
rect 883 200 887 204
rect 899 200 903 204
rect 42 -8 46 -4
rect 51 -8 55 -4
rect 60 -8 64 -4
rect 72 -8 76 -4
rect 81 -8 85 -4
rect 98 -8 102 -4
rect 107 -8 111 -4
rect 116 -8 120 -4
rect 128 -8 132 -4
rect 137 -8 141 -4
rect 154 -8 158 -4
rect 163 -8 167 -4
rect 172 -8 176 -4
rect 184 -8 188 -4
rect 193 -8 197 -4
rect 210 -8 214 -4
rect 219 -8 223 -4
rect 228 -8 232 -4
rect 240 -8 244 -4
rect 249 -8 253 -4
rect 266 -8 270 -4
rect 275 -8 279 -4
rect 284 -8 288 -4
rect 296 -8 300 -4
rect 305 -8 309 -4
rect 322 -8 326 -4
rect 331 -8 335 -4
rect 340 -8 344 -4
rect 352 -8 356 -4
rect 361 -8 365 -4
rect 378 -8 382 -4
rect 387 -8 391 -4
rect 396 -8 400 -4
rect 408 -8 412 -4
rect 417 -8 421 -4
rect 434 -8 438 -4
rect 443 -8 447 -4
rect 452 -8 456 -4
rect 464 -8 468 -4
rect 473 -8 477 -4
rect 490 -8 494 -4
rect 499 -8 503 -4
rect 508 -8 512 -4
rect 520 -8 524 -4
rect 529 -8 533 -4
rect 546 -8 550 -4
rect 555 -8 559 -4
rect 564 -8 568 -4
rect 576 -8 580 -4
rect 585 -8 589 -4
rect 602 -8 606 -4
rect 611 -8 615 -4
rect 620 -8 624 -4
rect 632 -8 636 -4
rect 641 -8 645 -4
rect 658 -8 662 -4
rect 667 -8 671 -4
rect 676 -8 680 -4
rect 688 -8 692 -4
rect 697 -8 701 -4
rect 714 -8 718 -4
rect 723 -8 727 -4
rect 732 -8 736 -4
rect 744 -8 748 -4
rect 753 -8 757 -4
rect 770 -8 774 -4
rect 779 -8 783 -4
rect 788 -8 792 -4
rect 800 -8 804 -4
rect 809 -8 813 -4
rect 826 -8 830 -4
rect 835 -8 839 -4
rect 844 -8 848 -4
rect 856 -8 860 -4
rect 865 -8 869 -4
<< polysilicon >>
rect 53 196 55 198
rect 74 196 76 198
rect 109 196 111 198
rect 130 196 132 198
rect 165 196 167 198
rect 186 196 188 198
rect 221 196 223 198
rect 242 196 244 198
rect 277 196 279 198
rect 298 196 300 198
rect 333 196 335 198
rect 354 196 356 198
rect 389 196 391 198
rect 410 196 412 198
rect 445 196 447 198
rect 466 196 468 198
rect 501 196 503 198
rect 522 196 524 198
rect 557 196 559 198
rect 578 196 580 198
rect 613 196 615 198
rect 634 196 636 198
rect 669 196 671 198
rect 690 196 692 198
rect 725 196 727 198
rect 746 196 748 198
rect 781 196 783 198
rect 802 196 804 198
rect 837 196 839 198
rect 858 196 860 198
rect 892 196 894 198
rect 900 196 902 198
rect 53 144 55 156
rect 74 144 76 156
rect 109 144 111 156
rect 130 144 132 156
rect 165 144 167 156
rect 186 144 188 156
rect 221 144 223 156
rect 242 144 244 156
rect 277 144 279 156
rect 298 144 300 156
rect 333 144 335 156
rect 354 144 356 156
rect 389 144 391 156
rect 410 144 412 156
rect 445 144 447 156
rect 466 144 468 156
rect 501 144 503 156
rect 522 144 524 156
rect 557 144 559 156
rect 578 144 580 156
rect 613 144 615 156
rect 634 144 636 156
rect 669 144 671 156
rect 690 144 692 156
rect 725 144 727 156
rect 746 144 748 156
rect 781 144 783 156
rect 802 144 804 156
rect 837 144 839 156
rect 858 144 860 156
rect 892 155 894 156
rect 900 155 902 156
rect 892 153 902 155
rect 53 140 63 144
rect 74 140 84 144
rect 109 140 119 144
rect 130 140 140 144
rect 165 140 175 144
rect 186 140 196 144
rect 221 140 231 144
rect 242 140 252 144
rect 277 140 287 144
rect 298 140 308 144
rect 333 140 343 144
rect 354 140 364 144
rect 389 140 399 144
rect 410 140 420 144
rect 445 140 455 144
rect 466 140 476 144
rect 501 140 511 144
rect 522 140 532 144
rect 557 140 567 144
rect 578 140 588 144
rect 613 140 623 144
rect 634 140 644 144
rect 669 140 679 144
rect 690 140 700 144
rect 725 140 735 144
rect 746 140 756 144
rect 781 140 791 144
rect 802 140 812 144
rect 837 140 847 144
rect 858 140 868 144
rect 48 128 50 131
rect 53 128 55 140
rect 69 128 71 131
rect 74 128 76 140
rect 104 128 106 131
rect 109 128 111 140
rect 125 128 127 131
rect 130 128 132 140
rect 160 128 162 131
rect 165 128 167 140
rect 181 128 183 131
rect 186 128 188 140
rect 216 128 218 131
rect 221 128 223 140
rect 237 128 239 131
rect 242 128 244 140
rect 272 128 274 131
rect 277 128 279 140
rect 293 128 295 131
rect 298 128 300 140
rect 328 128 330 131
rect 333 128 335 140
rect 349 128 351 131
rect 354 128 356 140
rect 384 128 386 131
rect 389 128 391 140
rect 405 128 407 131
rect 410 128 412 140
rect 440 128 442 131
rect 445 128 447 140
rect 461 128 463 131
rect 466 128 468 140
rect 496 128 498 131
rect 501 128 503 140
rect 517 128 519 131
rect 522 128 524 140
rect 552 128 554 131
rect 557 128 559 140
rect 573 128 575 131
rect 578 128 580 140
rect 608 128 610 131
rect 613 128 615 140
rect 629 128 631 131
rect 634 128 636 140
rect 664 128 666 131
rect 669 128 671 140
rect 685 128 687 131
rect 690 128 692 140
rect 720 128 722 131
rect 725 128 727 140
rect 741 128 743 131
rect 746 128 748 140
rect 776 128 778 131
rect 781 128 783 140
rect 797 128 799 131
rect 802 128 804 140
rect 832 128 834 131
rect 837 128 839 140
rect 853 128 855 131
rect 858 128 860 140
rect 892 135 894 153
rect 891 132 894 135
rect 891 131 902 132
rect 892 130 902 131
rect 892 128 894 130
rect 900 128 902 130
rect 48 106 50 108
rect 53 106 55 108
rect 69 106 71 108
rect 74 106 76 108
rect 104 106 106 108
rect 109 106 111 108
rect 125 106 127 108
rect 130 106 132 108
rect 160 106 162 108
rect 165 106 167 108
rect 181 106 183 108
rect 186 106 188 108
rect 216 106 218 108
rect 221 106 223 108
rect 237 106 239 108
rect 242 106 244 108
rect 272 106 274 108
rect 277 106 279 108
rect 293 106 295 108
rect 298 106 300 108
rect 328 106 330 108
rect 333 106 335 108
rect 349 106 351 108
rect 354 106 356 108
rect 384 106 386 108
rect 389 106 391 108
rect 405 106 407 108
rect 410 106 412 108
rect 440 106 442 108
rect 445 106 447 108
rect 461 106 463 108
rect 466 106 468 108
rect 496 106 498 108
rect 501 106 503 108
rect 517 106 519 108
rect 522 106 524 108
rect 552 106 554 108
rect 557 106 559 108
rect 573 106 575 108
rect 578 106 580 108
rect 608 106 610 108
rect 613 106 615 108
rect 629 106 631 108
rect 634 106 636 108
rect 664 106 666 108
rect 669 106 671 108
rect 685 106 687 108
rect 690 106 692 108
rect 720 106 722 108
rect 725 106 727 108
rect 741 106 743 108
rect 746 106 748 108
rect 776 106 778 108
rect 781 106 783 108
rect 797 106 799 108
rect 802 106 804 108
rect 832 106 834 108
rect 837 106 839 108
rect 853 106 855 108
rect 858 106 860 108
rect 892 106 894 108
rect 900 106 902 108
rect 48 88 50 90
rect 53 88 55 90
rect 69 88 71 90
rect 74 88 76 90
rect 104 88 106 90
rect 109 88 111 90
rect 125 88 127 90
rect 130 88 132 90
rect 160 88 162 90
rect 165 88 167 90
rect 181 88 183 90
rect 186 88 188 90
rect 216 88 218 90
rect 221 88 223 90
rect 237 88 239 90
rect 242 88 244 90
rect 272 88 274 90
rect 277 88 279 90
rect 293 88 295 90
rect 298 88 300 90
rect 328 88 330 90
rect 333 88 335 90
rect 349 88 351 90
rect 354 88 356 90
rect 384 88 386 90
rect 389 88 391 90
rect 405 88 407 90
rect 410 88 412 90
rect 440 88 442 90
rect 445 88 447 90
rect 461 88 463 90
rect 466 88 468 90
rect 496 88 498 90
rect 501 88 503 90
rect 517 88 519 90
rect 522 88 524 90
rect 552 88 554 90
rect 557 88 559 90
rect 573 88 575 90
rect 578 88 580 90
rect 608 88 610 90
rect 613 88 615 90
rect 629 88 631 90
rect 634 88 636 90
rect 664 88 666 90
rect 669 88 671 90
rect 685 88 687 90
rect 690 88 692 90
rect 720 88 722 90
rect 725 88 727 90
rect 741 88 743 90
rect 746 88 748 90
rect 776 88 778 90
rect 781 88 783 90
rect 797 88 799 90
rect 802 88 804 90
rect 832 88 834 90
rect 837 88 839 90
rect 853 88 855 90
rect 858 88 860 90
rect 48 65 50 68
rect 53 56 55 68
rect 69 65 71 68
rect 74 56 76 68
rect 104 65 106 68
rect 109 56 111 68
rect 125 65 127 68
rect 130 56 132 68
rect 160 65 162 68
rect 165 56 167 68
rect 181 65 183 68
rect 186 56 188 68
rect 216 65 218 68
rect 221 56 223 68
rect 237 65 239 68
rect 242 56 244 68
rect 272 65 274 68
rect 277 56 279 68
rect 293 65 295 68
rect 298 56 300 68
rect 328 65 330 68
rect 333 56 335 68
rect 349 65 351 68
rect 354 56 356 68
rect 384 65 386 68
rect 389 56 391 68
rect 405 65 407 68
rect 410 56 412 68
rect 440 65 442 68
rect 445 56 447 68
rect 461 65 463 68
rect 466 56 468 68
rect 496 65 498 68
rect 501 56 503 68
rect 517 65 519 68
rect 522 56 524 68
rect 552 65 554 68
rect 557 56 559 68
rect 573 65 575 68
rect 578 56 580 68
rect 608 65 610 68
rect 613 56 615 68
rect 629 65 631 68
rect 634 56 636 68
rect 664 65 666 68
rect 669 56 671 68
rect 685 65 687 68
rect 690 56 692 68
rect 720 65 722 68
rect 725 56 727 68
rect 741 65 743 68
rect 746 56 748 68
rect 776 65 778 68
rect 781 56 783 68
rect 797 65 799 68
rect 802 56 804 68
rect 832 65 834 68
rect 837 56 839 68
rect 853 65 855 68
rect 858 56 860 68
rect 53 52 63 56
rect 74 52 84 56
rect 109 52 119 56
rect 130 52 140 56
rect 165 52 175 56
rect 186 52 196 56
rect 221 52 231 56
rect 242 52 252 56
rect 277 52 287 56
rect 298 52 308 56
rect 333 52 343 56
rect 354 52 364 56
rect 389 52 399 56
rect 410 52 420 56
rect 445 52 455 56
rect 466 52 476 56
rect 501 52 511 56
rect 522 52 532 56
rect 557 52 567 56
rect 578 52 588 56
rect 613 52 623 56
rect 634 52 644 56
rect 669 52 679 56
rect 690 52 700 56
rect 725 52 735 56
rect 746 52 756 56
rect 781 52 791 56
rect 802 52 812 56
rect 837 52 847 56
rect 858 52 868 56
rect 53 40 55 52
rect 74 40 76 52
rect 109 40 111 52
rect 130 40 132 52
rect 165 40 167 52
rect 186 40 188 52
rect 221 40 223 52
rect 242 40 244 52
rect 277 40 279 52
rect 298 40 300 52
rect 333 40 335 52
rect 354 40 356 52
rect 389 40 391 52
rect 410 40 412 52
rect 445 40 447 52
rect 466 40 468 52
rect 501 40 503 52
rect 522 40 524 52
rect 557 40 559 52
rect 578 40 580 52
rect 613 40 615 52
rect 634 40 636 52
rect 669 40 671 52
rect 690 40 692 52
rect 725 40 727 52
rect 746 40 748 52
rect 781 40 783 52
rect 802 40 804 52
rect 837 40 839 52
rect 858 40 860 52
rect 53 -2 55 0
rect 74 -2 76 0
rect 109 -2 111 0
rect 130 -2 132 0
rect 165 -2 167 0
rect 186 -2 188 0
rect 221 -2 223 0
rect 242 -2 244 0
rect 277 -2 279 0
rect 298 -2 300 0
rect 333 -2 335 0
rect 354 -2 356 0
rect 389 -2 391 0
rect 410 -2 412 0
rect 445 -2 447 0
rect 466 -2 468 0
rect 501 -2 503 0
rect 522 -2 524 0
rect 557 -2 559 0
rect 578 -2 580 0
rect 613 -2 615 0
rect 634 -2 636 0
rect 669 -2 671 0
rect 690 -2 692 0
rect 725 -2 727 0
rect 746 -2 748 0
rect 781 -2 783 0
rect 802 -2 804 0
rect 837 -2 839 0
rect 858 -2 860 0
<< polycontact >>
rect 63 140 67 144
rect 84 140 88 144
rect 119 140 123 144
rect 140 140 144 144
rect 175 140 179 144
rect 196 140 200 144
rect 231 140 235 144
rect 252 140 256 144
rect 287 140 291 144
rect 308 140 312 144
rect 343 140 347 144
rect 364 140 368 144
rect 399 140 403 144
rect 420 140 424 144
rect 455 140 459 144
rect 476 140 480 144
rect 511 140 515 144
rect 532 140 536 144
rect 567 140 571 144
rect 588 140 592 144
rect 623 140 627 144
rect 644 140 648 144
rect 679 140 683 144
rect 700 140 704 144
rect 735 140 739 144
rect 756 140 760 144
rect 791 140 795 144
rect 812 140 816 144
rect 847 140 851 144
rect 868 140 872 144
rect 46 131 50 135
rect 67 131 71 135
rect 102 131 106 135
rect 123 131 127 135
rect 158 131 162 135
rect 179 131 183 135
rect 214 131 218 135
rect 235 131 239 135
rect 270 131 274 135
rect 291 131 295 135
rect 326 131 330 135
rect 347 131 351 135
rect 382 131 386 135
rect 403 131 407 135
rect 438 131 442 135
rect 459 131 463 135
rect 494 131 498 135
rect 515 131 519 135
rect 550 131 554 135
rect 571 131 575 135
rect 606 131 610 135
rect 627 131 631 135
rect 662 131 666 135
rect 683 131 687 135
rect 718 131 722 135
rect 739 131 743 135
rect 774 131 778 135
rect 795 131 799 135
rect 830 131 834 135
rect 851 131 855 135
rect 887 131 891 135
rect 46 61 50 65
rect 67 61 71 65
rect 102 61 106 65
rect 123 61 127 65
rect 158 61 162 65
rect 179 61 183 65
rect 214 61 218 65
rect 235 61 239 65
rect 270 61 274 65
rect 291 61 295 65
rect 326 61 330 65
rect 347 61 351 65
rect 382 61 386 65
rect 403 61 407 65
rect 438 61 442 65
rect 459 61 463 65
rect 494 61 498 65
rect 515 61 519 65
rect 550 61 554 65
rect 571 61 575 65
rect 606 61 610 65
rect 627 61 631 65
rect 662 61 666 65
rect 683 61 687 65
rect 718 61 722 65
rect 739 61 743 65
rect 774 61 778 65
rect 795 61 799 65
rect 830 61 834 65
rect 851 61 855 65
rect 63 52 67 56
rect 84 52 88 56
rect 119 52 123 56
rect 140 52 144 56
rect 175 52 179 56
rect 196 52 200 56
rect 231 52 235 56
rect 252 52 256 56
rect 287 52 291 56
rect 308 52 312 56
rect 343 52 347 56
rect 364 52 368 56
rect 399 52 403 56
rect 420 52 424 56
rect 455 52 459 56
rect 476 52 480 56
rect 511 52 515 56
rect 532 52 536 56
rect 567 52 571 56
rect 588 52 592 56
rect 623 52 627 56
rect 644 52 648 56
rect 679 52 683 56
rect 700 52 704 56
rect 735 52 739 56
rect 756 52 760 56
rect 791 52 795 56
rect 812 52 816 56
rect 847 52 851 56
rect 868 52 872 56
<< metal1 >>
rect 29 204 911 205
rect 29 200 42 204
rect 46 200 51 204
rect 55 200 60 204
rect 64 200 72 204
rect 76 200 81 204
rect 85 200 98 204
rect 102 200 107 204
rect 111 200 116 204
rect 120 200 128 204
rect 132 200 137 204
rect 141 200 154 204
rect 158 200 163 204
rect 167 200 172 204
rect 176 200 184 204
rect 188 200 193 204
rect 197 200 210 204
rect 214 200 219 204
rect 223 200 228 204
rect 232 200 240 204
rect 244 200 249 204
rect 253 200 266 204
rect 270 200 275 204
rect 279 200 284 204
rect 288 200 296 204
rect 300 200 305 204
rect 309 200 322 204
rect 326 200 331 204
rect 335 200 340 204
rect 344 200 352 204
rect 356 200 361 204
rect 365 200 378 204
rect 382 200 387 204
rect 391 200 396 204
rect 400 200 408 204
rect 412 200 417 204
rect 421 200 434 204
rect 438 200 443 204
rect 447 200 452 204
rect 456 200 464 204
rect 468 200 473 204
rect 477 200 490 204
rect 494 200 499 204
rect 503 200 508 204
rect 512 200 520 204
rect 524 200 529 204
rect 533 200 546 204
rect 550 200 555 204
rect 559 200 564 204
rect 568 200 576 204
rect 580 200 585 204
rect 589 200 602 204
rect 606 200 611 204
rect 615 200 620 204
rect 624 200 632 204
rect 636 200 641 204
rect 645 200 658 204
rect 662 200 667 204
rect 671 200 676 204
rect 680 200 688 204
rect 692 200 697 204
rect 701 200 714 204
rect 718 200 723 204
rect 727 200 732 204
rect 736 200 744 204
rect 748 200 753 204
rect 757 200 770 204
rect 774 200 779 204
rect 783 200 788 204
rect 792 200 800 204
rect 804 200 809 204
rect 813 200 826 204
rect 830 200 835 204
rect 839 200 844 204
rect 848 200 856 204
rect 860 200 865 204
rect 869 200 883 204
rect 887 200 899 204
rect 903 200 911 204
rect 29 199 911 200
rect 29 106 33 199
rect 48 196 52 199
rect 69 196 73 199
rect 104 196 108 199
rect 125 196 129 199
rect 160 196 164 199
rect 181 196 185 199
rect 216 196 220 199
rect 237 196 241 199
rect 272 196 276 199
rect 293 196 297 199
rect 328 196 332 199
rect 349 196 353 199
rect 384 196 388 199
rect 405 196 409 199
rect 440 196 444 199
rect 461 196 465 199
rect 496 196 500 199
rect 517 196 521 199
rect 552 196 556 199
rect 573 196 577 199
rect 608 196 612 199
rect 629 196 633 199
rect 664 196 668 199
rect 685 196 689 199
rect 720 196 724 199
rect 741 196 745 199
rect 776 196 780 199
rect 797 196 801 199
rect 832 196 836 199
rect 853 196 857 199
rect 887 196 891 199
rect 903 196 907 199
rect 56 144 60 156
rect 77 144 81 156
rect 112 144 116 156
rect 133 144 137 156
rect 168 144 172 156
rect 189 144 193 156
rect 224 144 228 156
rect 245 144 249 156
rect 280 144 284 156
rect 301 144 305 156
rect 336 144 340 156
rect 357 144 361 156
rect 392 144 396 156
rect 413 144 417 156
rect 448 144 452 156
rect 469 144 473 156
rect 504 144 508 156
rect 525 144 529 156
rect 560 144 564 156
rect 581 144 585 156
rect 616 144 620 156
rect 637 144 641 156
rect 672 144 676 156
rect 693 144 697 156
rect 728 144 732 156
rect 749 144 753 156
rect 784 144 788 156
rect 805 144 809 156
rect 840 144 844 156
rect 861 144 865 156
rect 36 140 60 144
rect 67 140 81 144
rect 88 140 116 144
rect 123 140 137 144
rect 144 140 172 144
rect 179 140 193 144
rect 200 140 228 144
rect 235 140 249 144
rect 256 140 284 144
rect 291 140 305 144
rect 312 140 340 144
rect 347 140 361 144
rect 368 140 396 144
rect 403 140 417 144
rect 424 140 452 144
rect 459 140 473 144
rect 480 140 508 144
rect 515 140 529 144
rect 536 140 564 144
rect 571 140 585 144
rect 592 140 620 144
rect 627 140 641 144
rect 648 140 676 144
rect 683 140 697 144
rect 704 140 732 144
rect 739 140 753 144
rect 760 140 788 144
rect 795 140 809 144
rect 816 140 844 144
rect 851 140 865 144
rect 36 106 40 140
rect 50 131 51 135
rect 56 128 60 140
rect 71 131 72 135
rect 77 128 81 140
rect 106 131 107 135
rect 112 128 116 140
rect 127 131 128 135
rect 133 128 137 140
rect 162 131 163 135
rect 168 128 172 140
rect 183 131 184 135
rect 189 128 193 140
rect 218 131 219 135
rect 224 128 228 140
rect 239 131 240 135
rect 245 128 249 140
rect 274 131 275 135
rect 280 128 284 140
rect 295 131 296 135
rect 301 128 305 140
rect 330 131 331 135
rect 336 128 340 140
rect 351 131 352 135
rect 357 128 361 140
rect 386 131 387 135
rect 392 128 396 140
rect 407 131 408 135
rect 413 128 417 140
rect 442 131 443 135
rect 448 128 452 140
rect 463 131 464 135
rect 469 128 473 140
rect 498 131 499 135
rect 504 128 508 140
rect 519 131 520 135
rect 525 128 529 140
rect 554 131 555 135
rect 560 128 564 140
rect 575 131 576 135
rect 581 128 585 140
rect 610 131 611 135
rect 616 128 620 140
rect 631 131 632 135
rect 637 128 641 140
rect 666 131 667 135
rect 672 128 676 140
rect 687 131 688 135
rect 693 128 697 140
rect 722 131 723 135
rect 728 128 732 140
rect 743 131 744 135
rect 749 128 753 140
rect 778 131 779 135
rect 784 128 788 140
rect 799 131 800 135
rect 805 128 809 140
rect 834 131 835 135
rect 840 128 844 140
rect 850 131 851 135
rect 861 128 865 140
rect 868 136 891 140
rect 887 135 891 136
rect 895 135 899 156
rect 895 131 913 135
rect 895 128 899 131
rect 29 92 40 106
rect 29 -3 33 92
rect 36 56 40 92
rect 43 105 47 108
rect 64 105 68 108
rect 99 105 103 108
rect 120 105 124 108
rect 155 105 159 108
rect 176 105 180 108
rect 211 105 215 108
rect 232 105 236 108
rect 267 105 271 108
rect 288 105 292 108
rect 323 105 327 108
rect 344 105 348 108
rect 379 105 383 108
rect 400 105 404 108
rect 435 105 439 108
rect 456 105 460 108
rect 491 105 495 108
rect 512 105 516 108
rect 547 105 551 108
rect 568 105 572 108
rect 603 105 607 108
rect 624 105 628 108
rect 659 105 663 108
rect 680 105 684 108
rect 715 105 719 108
rect 736 105 740 108
rect 771 105 775 108
rect 792 105 796 108
rect 827 105 831 108
rect 848 105 852 108
rect 887 105 891 108
rect 903 105 907 108
rect 43 104 912 105
rect 43 100 51 104
rect 55 100 60 104
rect 64 100 72 104
rect 76 100 81 104
rect 85 100 98 104
rect 102 100 107 104
rect 111 100 116 104
rect 120 100 128 104
rect 132 100 137 104
rect 141 100 154 104
rect 158 100 163 104
rect 167 100 172 104
rect 176 100 184 104
rect 188 100 193 104
rect 197 100 210 104
rect 214 100 219 104
rect 223 100 228 104
rect 232 100 240 104
rect 244 100 249 104
rect 253 100 266 104
rect 270 100 275 104
rect 279 100 284 104
rect 288 100 296 104
rect 300 100 305 104
rect 309 100 322 104
rect 326 100 331 104
rect 335 100 340 104
rect 344 100 352 104
rect 356 100 361 104
rect 365 100 378 104
rect 382 100 387 104
rect 391 100 396 104
rect 400 100 408 104
rect 412 100 417 104
rect 421 100 434 104
rect 438 100 443 104
rect 447 100 452 104
rect 456 100 464 104
rect 468 100 473 104
rect 477 100 490 104
rect 494 100 499 104
rect 503 100 508 104
rect 512 100 520 104
rect 524 100 529 104
rect 533 100 546 104
rect 550 100 555 104
rect 559 100 564 104
rect 568 100 576 104
rect 580 100 585 104
rect 589 100 602 104
rect 606 100 611 104
rect 615 100 620 104
rect 624 100 632 104
rect 636 100 641 104
rect 645 100 658 104
rect 662 100 667 104
rect 671 100 676 104
rect 680 100 688 104
rect 692 100 697 104
rect 701 100 714 104
rect 718 100 723 104
rect 727 100 732 104
rect 736 100 744 104
rect 748 100 753 104
rect 757 100 770 104
rect 774 100 779 104
rect 783 100 788 104
rect 792 100 800 104
rect 804 100 809 104
rect 813 100 826 104
rect 830 100 835 104
rect 839 100 844 104
rect 848 100 856 104
rect 860 100 868 104
rect 872 100 883 104
rect 887 100 899 104
rect 903 100 912 104
rect 43 96 912 100
rect 43 92 51 96
rect 55 92 60 96
rect 64 92 72 96
rect 76 92 81 96
rect 85 92 98 96
rect 102 92 107 96
rect 111 92 116 96
rect 120 92 128 96
rect 132 92 137 96
rect 141 92 154 96
rect 158 92 163 96
rect 167 92 172 96
rect 176 92 184 96
rect 188 92 193 96
rect 197 92 210 96
rect 214 92 219 96
rect 223 92 228 96
rect 232 92 240 96
rect 244 92 249 96
rect 253 92 266 96
rect 270 92 275 96
rect 279 92 284 96
rect 288 92 296 96
rect 300 92 305 96
rect 309 92 322 96
rect 326 92 331 96
rect 335 92 340 96
rect 344 92 352 96
rect 356 92 361 96
rect 365 92 378 96
rect 382 92 387 96
rect 391 92 396 96
rect 400 92 408 96
rect 412 92 417 96
rect 421 92 434 96
rect 438 92 443 96
rect 447 92 452 96
rect 456 92 464 96
rect 468 92 473 96
rect 477 92 490 96
rect 494 92 499 96
rect 503 92 508 96
rect 512 92 520 96
rect 524 92 529 96
rect 533 92 546 96
rect 550 92 555 96
rect 559 92 564 96
rect 568 92 576 96
rect 580 92 585 96
rect 589 92 602 96
rect 606 92 611 96
rect 615 92 620 96
rect 624 92 632 96
rect 636 92 641 96
rect 645 92 658 96
rect 662 92 667 96
rect 671 92 676 96
rect 680 92 688 96
rect 692 92 697 96
rect 701 92 714 96
rect 718 92 723 96
rect 727 92 732 96
rect 736 92 744 96
rect 748 92 753 96
rect 757 92 770 96
rect 774 92 779 96
rect 783 92 788 96
rect 792 92 800 96
rect 804 92 809 96
rect 813 92 826 96
rect 830 92 835 96
rect 839 92 844 96
rect 848 92 856 96
rect 860 92 868 96
rect 872 92 883 96
rect 887 92 899 96
rect 903 92 912 96
rect 43 91 912 92
rect 43 88 47 91
rect 64 88 68 91
rect 99 88 103 91
rect 120 88 124 91
rect 155 88 159 91
rect 176 88 180 91
rect 211 88 215 91
rect 232 88 236 91
rect 267 88 271 91
rect 288 88 292 91
rect 323 88 327 91
rect 344 88 348 91
rect 379 88 383 91
rect 400 88 404 91
rect 435 88 439 91
rect 456 88 460 91
rect 491 88 495 91
rect 512 88 516 91
rect 547 88 551 91
rect 568 88 572 91
rect 603 88 607 91
rect 624 88 628 91
rect 659 88 663 91
rect 680 88 684 91
rect 715 88 719 91
rect 736 88 740 91
rect 771 88 775 91
rect 792 88 796 91
rect 827 88 831 91
rect 848 88 852 91
rect 50 61 51 65
rect 56 56 60 68
rect 71 61 72 65
rect 77 56 81 68
rect 106 61 107 65
rect 112 56 116 68
rect 127 61 128 65
rect 133 56 137 68
rect 162 61 163 65
rect 168 56 172 68
rect 183 61 184 65
rect 189 56 193 68
rect 218 61 219 65
rect 224 56 228 68
rect 239 61 240 65
rect 245 56 249 68
rect 274 61 275 65
rect 280 56 284 68
rect 295 61 296 65
rect 301 56 305 68
rect 330 61 331 65
rect 336 56 340 68
rect 351 61 352 65
rect 357 56 361 68
rect 386 61 387 65
rect 392 56 396 68
rect 407 61 408 65
rect 413 56 417 68
rect 442 61 443 65
rect 448 56 452 68
rect 463 61 464 65
rect 469 56 473 68
rect 498 61 499 65
rect 504 56 508 68
rect 519 61 520 65
rect 525 56 529 68
rect 554 61 555 65
rect 560 56 564 68
rect 575 61 576 65
rect 581 56 585 68
rect 610 61 611 65
rect 616 56 620 68
rect 631 61 632 65
rect 637 56 641 68
rect 666 61 667 65
rect 672 56 676 68
rect 687 61 688 65
rect 693 56 697 68
rect 722 61 723 65
rect 728 56 732 68
rect 743 61 744 65
rect 749 56 753 68
rect 778 61 779 65
rect 784 56 788 68
rect 799 61 800 65
rect 805 56 809 68
rect 834 61 835 65
rect 840 56 844 68
rect 850 61 851 65
rect 861 56 865 68
rect 36 52 60 56
rect 67 52 81 56
rect 88 52 116 56
rect 123 52 137 56
rect 144 52 172 56
rect 179 52 193 56
rect 200 52 228 56
rect 235 52 249 56
rect 256 52 284 56
rect 291 52 305 56
rect 312 52 340 56
rect 347 52 361 56
rect 368 52 396 56
rect 403 52 417 56
rect 424 52 452 56
rect 459 52 473 56
rect 480 52 508 56
rect 515 52 529 56
rect 536 52 564 56
rect 571 52 585 56
rect 592 52 620 56
rect 627 52 641 56
rect 648 52 676 56
rect 683 52 697 56
rect 704 52 732 56
rect 739 52 753 56
rect 760 52 788 56
rect 795 52 809 56
rect 816 52 844 56
rect 851 52 865 56
rect 868 56 872 60
rect 56 40 60 52
rect 77 40 81 52
rect 112 40 116 52
rect 133 40 137 52
rect 168 40 172 52
rect 189 40 193 52
rect 224 40 228 52
rect 245 40 249 52
rect 280 40 284 52
rect 301 40 305 52
rect 336 40 340 52
rect 357 40 361 52
rect 392 40 396 52
rect 413 40 417 52
rect 448 40 452 52
rect 469 40 473 52
rect 504 40 508 52
rect 525 40 529 52
rect 560 40 564 52
rect 581 40 585 52
rect 616 40 620 52
rect 637 40 641 52
rect 672 40 676 52
rect 693 40 697 52
rect 728 40 732 52
rect 749 40 753 52
rect 784 40 788 52
rect 805 40 809 52
rect 840 40 844 52
rect 861 40 865 52
rect 48 -3 52 0
rect 69 -3 73 0
rect 104 -3 108 0
rect 125 -3 129 0
rect 160 -3 164 0
rect 181 -3 185 0
rect 216 -3 220 0
rect 237 -3 241 0
rect 272 -3 276 0
rect 293 -3 297 0
rect 328 -3 332 0
rect 349 -3 353 0
rect 384 -3 388 0
rect 405 -3 409 0
rect 440 -3 444 0
rect 461 -3 465 0
rect 496 -3 500 0
rect 517 -3 521 0
rect 552 -3 556 0
rect 573 -3 577 0
rect 608 -3 612 0
rect 629 -3 633 0
rect 664 -3 668 0
rect 685 -3 689 0
rect 720 -3 724 0
rect 741 -3 745 0
rect 776 -3 780 0
rect 797 -3 801 0
rect 832 -3 836 0
rect 853 -3 857 0
rect 29 -4 876 -3
rect 29 -8 42 -4
rect 46 -8 51 -4
rect 55 -8 60 -4
rect 64 -8 72 -4
rect 76 -8 81 -4
rect 85 -8 98 -4
rect 102 -8 107 -4
rect 111 -8 116 -4
rect 120 -8 128 -4
rect 132 -8 137 -4
rect 141 -8 154 -4
rect 158 -8 163 -4
rect 167 -8 172 -4
rect 176 -8 184 -4
rect 188 -8 193 -4
rect 197 -8 210 -4
rect 214 -8 219 -4
rect 223 -8 228 -4
rect 232 -8 240 -4
rect 244 -8 249 -4
rect 253 -8 266 -4
rect 270 -8 275 -4
rect 279 -8 284 -4
rect 288 -8 296 -4
rect 300 -8 305 -4
rect 309 -8 322 -4
rect 326 -8 331 -4
rect 335 -8 340 -4
rect 344 -8 352 -4
rect 356 -8 361 -4
rect 365 -8 378 -4
rect 382 -8 387 -4
rect 391 -8 396 -4
rect 400 -8 408 -4
rect 412 -8 417 -4
rect 421 -8 434 -4
rect 438 -8 443 -4
rect 447 -8 452 -4
rect 456 -8 464 -4
rect 468 -8 473 -4
rect 477 -8 490 -4
rect 494 -8 499 -4
rect 503 -8 508 -4
rect 512 -8 520 -4
rect 524 -8 529 -4
rect 533 -8 546 -4
rect 550 -8 555 -4
rect 559 -8 564 -4
rect 568 -8 576 -4
rect 580 -8 585 -4
rect 589 -8 602 -4
rect 606 -8 611 -4
rect 615 -8 620 -4
rect 624 -8 632 -4
rect 636 -8 641 -4
rect 645 -8 658 -4
rect 662 -8 667 -4
rect 671 -8 676 -4
rect 680 -8 688 -4
rect 692 -8 697 -4
rect 701 -8 714 -4
rect 718 -8 723 -4
rect 727 -8 732 -4
rect 736 -8 744 -4
rect 748 -8 753 -4
rect 757 -8 770 -4
rect 774 -8 779 -4
rect 783 -8 788 -4
rect 792 -8 800 -4
rect 804 -8 809 -4
rect 813 -8 826 -4
rect 830 -8 835 -4
rect 839 -8 844 -4
rect 848 -8 856 -4
rect 860 -8 865 -4
rect 869 -8 876 -4
rect 29 -9 876 -8
<< m2contact >>
rect 46 131 50 135
rect 67 131 71 135
rect 102 131 106 135
rect 123 131 127 135
rect 158 131 162 135
rect 179 131 183 135
rect 214 131 218 135
rect 235 131 239 135
rect 270 131 274 135
rect 291 131 295 135
rect 326 131 330 135
rect 347 131 351 135
rect 382 131 386 135
rect 403 131 407 135
rect 438 131 442 135
rect 459 131 463 135
rect 494 131 498 135
rect 515 131 519 135
rect 550 131 554 135
rect 571 131 575 135
rect 606 131 610 135
rect 627 131 631 135
rect 662 131 666 135
rect 683 131 687 135
rect 718 131 722 135
rect 739 131 743 135
rect 774 131 778 135
rect 795 131 799 135
rect 830 131 834 135
rect 851 131 855 135
rect 868 140 872 144
rect 46 61 50 65
rect 67 61 71 65
rect 102 61 106 65
rect 123 61 127 65
rect 158 61 162 65
rect 179 61 183 65
rect 214 61 218 65
rect 235 61 239 65
rect 270 61 274 65
rect 291 61 295 65
rect 326 61 330 65
rect 347 61 351 65
rect 382 61 386 65
rect 403 61 407 65
rect 438 61 442 65
rect 459 61 463 65
rect 494 61 498 65
rect 515 61 519 65
rect 550 61 554 65
rect 571 61 575 65
rect 606 61 610 65
rect 627 61 631 65
rect 662 61 666 65
rect 683 61 687 65
rect 718 61 722 65
rect 739 61 743 65
rect 774 61 778 65
rect 795 61 799 65
rect 830 61 834 65
rect 851 61 855 65
rect 868 52 872 56
<< metal2 >>
rect 36 131 46 135
rect 50 131 67 135
rect 71 131 102 135
rect 106 131 123 135
rect 127 131 158 135
rect 162 131 179 135
rect 183 131 214 135
rect 218 131 235 135
rect 239 131 270 135
rect 274 131 291 135
rect 295 131 326 135
rect 330 131 347 135
rect 351 131 382 135
rect 386 131 403 135
rect 407 131 438 135
rect 442 131 459 135
rect 463 131 494 135
rect 498 131 515 135
rect 519 131 550 135
rect 554 131 571 135
rect 575 131 606 135
rect 610 131 627 135
rect 631 131 662 135
rect 666 131 683 135
rect 687 131 718 135
rect 722 131 739 135
rect 743 131 774 135
rect 778 131 795 135
rect 799 131 830 135
rect 834 131 851 135
rect 36 106 40 131
rect 29 92 40 106
rect 36 65 40 92
rect 36 61 46 65
rect 50 61 67 65
rect 71 61 102 65
rect 106 61 123 65
rect 127 61 158 65
rect 162 61 179 65
rect 183 61 214 65
rect 218 61 235 65
rect 239 61 270 65
rect 274 61 291 65
rect 295 61 326 65
rect 330 61 347 65
rect 351 61 382 65
rect 386 61 403 65
rect 407 61 438 65
rect 442 61 459 65
rect 463 61 494 65
rect 498 61 515 65
rect 519 61 550 65
rect 554 61 571 65
rect 575 61 606 65
rect 610 61 627 65
rect 631 61 662 65
rect 666 61 683 65
rect 687 61 718 65
rect 722 61 739 65
rect 743 61 774 65
rect 778 61 795 65
rect 799 61 830 65
rect 834 61 851 65
rect 868 56 872 140
<< m1p >>
rect 895 145 899 149
rect 868 136 891 140
rect 887 135 891 136
<< labels >>
rlabel metal1 38 202 38 202 5 vdd!
rlabel metal2 29 92 29 106 3 vcoctrl
rlabel metal1 859 98 859 98 1 gnd!
rlabel metal1 913 131 913 135 7 fout
<< end >>
